

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.all;
USE ieee.numeric_std.ALL;

entity VideoGame is

      Port (Clickbuttons : in STD_LOGIC_VECTOR (4 downto 0);
            display, Halfclock : in std_logic;
            pokemonFramer: in std_logic_vector(8 downto 0);
            Rin, Bin, Gin : out std_logic_vector(3 downto 0);
            Pokemonchooser : in std_logic_vector(3 downto 0);
            T1P1: in std_logic_vector(8 downto 0);
            T1P2: in std_logic_vector(8 downto 0);
            T2P1: in std_logic_vector(8 downto 0);
            T2P2: in std_logic_vector(8 downto 0);
            ssingle : in std_logic;
            Angriff : in std_logic_vector (2 downto 0);
            Ddamage : in std_logic;
            Pokemonnumbers : in std_logic_vector(2 downto 0);
            Sschaden : in std_logic_vector(4 downto 0);
            Winner : in std_logic;
            PAliveStatus : in std_logic_vector(3 downto 0);
            PokemonStats : in std_logic_vector(19 downto 0);
            menu : in STD_LOGIC_VECTOR (2 downto 0);
            Bmenu : in STD_LOGIC_VECTOR (2 downto 0);
            pixel_X : in std_logic_vector(10 downto 0);
            pixel_Y : in std_logic_vector(9 downto 0));

end VideoGame;

architecture Behavioral of VideoGame is

signal TeamOne: std_logic_vector(2 downto 0);

type Feuer is array (0 to 12, 0 to 33) of std_logic_vector(5 downto 0);
type Wasser is array (0 to 44, 0 to 19) of std_logic_vector(5 downto 0);
type Pflanze is array (0 to 22, 0 to 26) of std_logic_vector(5 downto 0);
type Normale is array (0 to 16, 0 to 19) of std_logic_vector(5 downto 0);
type wins is array (0 to 33, 0 to 90) of std_logic;
type plays is array(0 to 38, 0 to 88) of std_logic;
type team is array(0 to 33, 0 to 87) of std_logic;
type s1 is array(0 to 33, 0 to 15) of std_logic;
type s2 is array(0 to 33, 0 to 22) of std_logic;
type choose is array(0 to 37, 0 to 111) of std_logic;
type PokemonBits is array (0 to 159, 0 to 281) of std_logic_vector(5 downto 0);
type Hp is array (0 to 56, 0 to 62) of std_logic_vector(5 downto 0);
type At is array (0 to 51, 0 to 70) of std_logic_vector(5 downto 0);
type Def is array (0 to 44, 0 to 81) of std_logic_vector(5 downto 0);
type Sp is array (0 to 54, 0 to 62) of std_logic_vector(5 downto 0);
type MegaPunch is array (0 to 28, 0 to 136) of std_logic;
type FireBlast is array (0 to 24, 0 to 96) of std_logic;
type LeafBlade is array (0 to 24, 0 to 115) of std_logic;
type Surf is array (0 to 22, 0 to 47) of std_logic;
type Nott is array (0 to 16, 0 to 36) of std_logic;
type VeryEffective is array (0 to 21, 0 to 155) of std_logic;
type SinglePlayer is array (0 to 26, 0 to 131) of std_logic;
type Multiplayer is array (0 to 26, 0 to 124) of std_logic;

type Pokemon is array (0 to 55, 0 to 55) of std_logic_vector(5 downto 0);


constant pflanzeString : pflanze:= (("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","011100","011100","000100","000100","000100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","011100","000100","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000100","000100","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","011100","011100","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","000100","000100","000100","011100","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","000100","011100","011100","011100","011100","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000100","000100","011100","011100","011100","011100","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","011100","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","011100","011100","000100","000100","000100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","011100","000100","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000100","000100","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"));

constant wasserString : wasser:= (("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","101111","101111","101111","000000","000000","000000","000000","101111","101111","101111","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","101111","101111","000000","000000","101111","101111","000000","000000","111111","000000"),
("000000","000000","000000","000000","000000","000000","000000","101111","111111","011011","000111","000111","011011","011011","000111","000111","011011","111111","101111","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","001011","000111","000111","000111","000111","000111","000111","000111","000111","001011","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","101011","000111","001011","001011","001011","001011","001011","001011","001011","001011","000111","101011","000000"),
("000000","000000","000000","000000","000000","000000","000000","001011","000111","000111","001011","001011","000111","000111","001011","001011","000111","000111","001011","000000"),
("000000","000000","000000","000000","000000","000000","000000","001011","001011","000111","000111","001011","000111","000111","001011","000111","000111","001011","001011","000000"),
("000000","000000","000000","000000","000000","000000","000000","001011","001011","011011","001011","011011","011011","011011","011011","001011","011011","001011","001011","000000"),
("000000","000000","000000","000000","000000","000000","000000","101111","000111","001011","001011","000111","001011","001011","000111","001011","001011","000111","011011","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000110","000111","101111","011011","000111","000111","011011","101111","001011","011011","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001011","000111","000111","000111","000111","001011","101011","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001011","001011","001011","001011","001011","000111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","001011","001011","001011","001011","000111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000111","000111","000111","000111","000111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","001011","001011","001011","001011","001011","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001011","001011","001011","001011","001011","000111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000111","000111","000111","000111","000111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","001011","001011","001011","001011","001011","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","001011","001011","001011","001011","000111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001011","000111","000111","000111","000111","001011","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001011","001011","001011","001011","001011","001011","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","001011","001011","001011","001011","000111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000111","000111","000111","000111","001011","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001011","001011","001011","001011","001011","001011","000000","000000","000000","000000"),
("000000","000000","101111","101111","101111","000000","000000","000000","000000","101011","000111","001011","001011","001011","001011","000111","000000","000000","000000","000000"),
("000000","111111","000000","000000","101111","101111","000000","000000","101111","101111","000111","000111","000111","000111","000111","001011","000000","000000","000000","000000"),
("000000","101111","111111","011011","000111","000111","011011","011011","000111","000111","000111","001011","001011","001011","001011","000111","000000","000000","000000","000000"),
("000000","000000","001011","000111","000111","000111","000111","000111","000111","000111","000111","001011","000111","001011","001011","000111","000000","000000","000000","000000"),
("000000","101011","000111","001011","001011","001011","001011","001011","001011","001011","001011","001011","000111","000111","000111","000111","000000","000000","000000","000000"),
("000000","001011","000111","000111","001011","001011","000111","000111","001011","001011","000111","000111","000111","001011","001011","000111","000000","000000","000000","000000"),
("000000","001011","001011","000111","000111","001011","000111","000111","001011","000111","000111","001011","000111","001011","001011","000111","000000","000000","000000","000000"),
("000000","001011","001011","011011","001011","011011","011011","011011","011011","001011","011011","001011","000111","000111","000111","000111","000000","000000","000000","000000"),
("000000","011011","000111","001011","001011","000111","001011","001011","000111","001011","001011","000111","001011","001011","001011","000111","000000","000000","000000","000000"),
("000000","000000","011011","000111","101111","011011","000111","000111","011011","101111","000111","000111","001011","001011","001011","000111","000000","000000","000000","000000"),
("000000","000000","000000","000000","001011","000111","000111","000111","000111","001011","000111","000111","000111","000111","000111","000111","000000","000000","000000","000000"),
("000000","000000","000000","000000","001011","001011","001011","001011","001011","000111","000111","001011","001011","001011","001011","000111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000111","001011","001011","001011","001011","000111","000111","001011","001011","001011","001011","000111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000000","000000","000000","000000"),
("000000","000000","000000","000000","001011","001011","001011","001011","001011","000111","000111","001011","001011","001011","001011","001011","000000","000000","000000","000000"),
("000000","000000","000000","000000","001011","011011","001011","001011","011011","000111","000111","011011","001011","001011","011011","001011","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"));

constant feuerString : feuer:= (("000000","110000","110000","000000","000000","000000","000000","110000","111100","110000","111100","000000","000000","000000","000000","111100","000000","000000","000000","111100","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("110000","111100","000000","000000","110000","111100","110000","111100","110000","000000","000000","000000","111100","110000","111100","000000","000000","000000","111100","110000","111100","110000","000000","000000","000000","000000","111100","110000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","111100","110000","110000","110000","111100","111100","111100","110000","110000","000000","000000","000000","000000","111100","110000","111100","110000","111100","110000","000000","000000","111100","110000","111111","110000","000000","000000","000000","000000","000000"),
("000000","000000","111100","000000","110000","110000","110000","111100","111100","110000","110000","111100","000000","000000","000000","000000","000000","110000","111100","110000","111100","110000","110000","110000","111100","110000","110000","110000","000000","110000","000000","000000","000000","000000"),
("000000","000000","000000","110000","110000","110000","110000","110000","110000","110000","110000","110000","000000","000000","000000","000000","000000","110000","111100","111100","110000","110000","110000","110000","110000","110000","110000","000000","000000","000000","000000","000000","000000","000000"),
("000000","110000","000000","110000","000000","110000","110000","110000","110000","110000","000000","111100","110000","110000","110000","000000","110000","111100","111100","110000","110000","111100","110000","110000","110000","110000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","110000","000000","000000","110000","111100","110000","111100","110000","110000","110000","110000","111100","110000","111100","111100","111100","111100","110000","110000","111100","000000","111100","110000","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("110000","110000","111100","110000","111100","110000","111100","110000","111100","000000","110000","110000","110000","111100","111100","111100","111100","110000","111100","110000","000000","000000","000000","000000","000000","000000","000000","110000","110000","110000","000000","000000","000000","000000"),
("110000","111100","110000","111100","110000","111100","111100","111100","111100","111100","000000","110000","110000","110000","111100","111100","111100","111100","110000","110000","110000","111100","000000","000000","000000","110000","111100","111100","111100","111100","110000","110000","110000","000000"),
("111100","110000","111100","110000","111100","110000","111100","111100","111100","111100","111100","111100","110000","111100","110000","111100","110000","110000","110000","110000","110000","111100","000000","110000","110000","111100","111100","111100","111100","111100","111100","111100","111100","110000"),
("110000","110000","110000","111100","110000","111100","110000","111100","110000","111100","111100","111100","111100","110000","111100","110000","110000","110000","000000","110000","111100","000000","110000","111100","111100","111100","111100","111100","110000","111100","110000","111100","110000","111100"),
("110000","110000","110000","110000","110000","110000","110000","110000","111100","110000","111100","111100","110000","111100","110000","110000","110000","000000","000000","000000","000000","000000","110000","111100","111100","111100","111100","110000","111100","110000","111100","110000","111100","110000"),
("110000","110000","110000","110000","110000","110000","110000","110000","110000","111100","111100","110000","111100","110000","111100","110000","110000","000000","000000","000000","000000","000000","110000","111100","111100","111100","110000","111100","110000","110000","110000","110000","110000","110000"));

constant normaleString : normale:= (("101001","101010","101010","010101","000000","000000","000000","000000","101010","111111","111111","111111","101010","111111","111111","111111","111111","101010","000000","000000"),
("101010","101010","111111","101010","101010","101010","010101","101010","111111","111111","111111","111111","101010","111111","111111","101010","101010","111111","111111","000000"),
("000000","010101","101011","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","101010","111111","000000"),
("000000","000000","101010","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","101010","000000","000000"),
("000000","000000","101001","111111","111111","010101","010101","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","101010","000000","000000"),
("000000","000000","010101","111111","111111","010101","010101","111111","010101","010101","111111","000000","010101","111111","111111","111111","111111","010101","000000","000000"),
("010101","101010","101010","111111","111111","010101","010101","111111","010101","010101","111111","010101","010101","111111","010101","101010","111111","101010","101010","000000"),
("010101","101010","111111","111111","111111","010101","010101","111111","010101","010101","111111","010101","010101","111111","010101","101010","111111","111111","111010","000000"),
("111111","111111","111111","111111","111111","010101","010101","111111","010101","010101","111111","010101","010101","111111","010101","101010","111111","111111","111111","111111"),
("111111","111111","111111","111111","111111","010101","010101","101010","010101","010101","101010","010101","010101","111111","010101","101010","111111","111111","111111","111111"),
("010101","101010","111111","111111","111111","010101","010101","010101","010101","010101","101010","010101","010101","010101","101010","111111","111111","111111","101010","010101"),
("101010","010101","101010","111111","111111","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","111111","111111","101010","111111","000000"),
("000000","101010","010101","111111","111111","010101","010101","000000","010101","010101","010101","010101","010101","000000","101010","111111","111111","010101","000000","000000"),
("000000","000000","101010","111111","111111","111111","111111","010101","010101","010101","010101","010101","000000","101010","111111","111111","111111","101010","000000","000000"),
("000000","000000","101010","111111","111111","111111","111111","111111","010101","010101","010101","010101","101010","111111","111111","111111","111111","101010","000000","000000"),
("000000","111111","101010","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","101010","111111","000000"),
("000000","101010","111111","101010","101010","010101","010101","101010","111111","111111","111111","111111","101010","010101","000000","000000","000000","000000","000000","000000"));


constant teamString : team:= (('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','1','1','0','0','0','0','0','0','1','1','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','1','0','0','0','0','0','0','1','1','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','1','1','1','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','1','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0'),
('0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0'),
('0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','0','0','1','1','1','1','1','1','1','0','1','1','1','1','1','1','1','1','0','1','1','1','1','1','1','1','1','0','1','1','1','1','1','1','1','1','0'),
('0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','1','1','1','1','1','1','1','0','0','0','1','1','0','0','0','0','0','0','1','1','1','1','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0'),
('0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0'),
('0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0'),
('0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','1','1','1','1','1','1','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','0'),
('0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','0','0','1','1','1','0','0','1','1','1','1','1','1','0','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','0'),
('0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0'),
('0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','0','1','1','1','1','1','1','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','0','1','1','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));


constant playsString : plays := (('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','1','1','1','1','1','1','1','1','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0'),
('0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0'),
('0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','0','0','1','1','1','1','1','1','1','0','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','1','1','0','0','0','0','1','1','1','1','1','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','1','1','1','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','1','1','0','0','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','1','1','1','0','0','1','1','1','1','1','1','0','0','1','1','1','1','1','1','0','0'),
('0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0'),
('0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0'),
('0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','0','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','1','1','1'),
('0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','1','1'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','1','0'),
('0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','0','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','1','0'),
('1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','1','1','1','1','1','1','1','1','1','0','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','0','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0'),
('1','1','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','0','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0'),
('0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));


constant winsString : wins := (('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','1','1','1','1','1','1','1','0','1','1','1','0','0','0','0','1','1','1','1','1','1','1','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','1','1','1','1','1','1','1','0','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0'),
('0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0','1','1','1','1','1','1','0','0','0','0'),
('0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','1','1','1','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0'),
('0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','1','0','0','0'),
('0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','1','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','1','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','1','1','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0'),
('0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));

constant oneString : s1:= (('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0'),
('0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0'),
('0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0'),
('0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0'),
('0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0'),
('0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));


constant twoString : s2:= (('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0'),
('0','0','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0'),
('0','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0'),
('0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0'),
('0','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));

constant chooseString : choose:= (('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','1','1','0','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','1','1','1','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
('0','0','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0'),
('0','1','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0'),
('0','1','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0'),
('0','1','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1'),
('0','1','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','1','1','0','1','1','1','1','1','1'),
('0','1','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','1','1','1','0','0','1','1','1','1','1'),
('0','1','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','1','0','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','0'),
('0','1','1','1','1','1','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','1','0','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','1','1','1','1','1','1','0','0','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','1','1','1','0','0','0'),
('0','1','1','1','1','1','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','0','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0'),
('0','1','1','1','1','1','1','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0'),
('0','1','1','1','1','1','1','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','1','1','1','1','1','0','0','0','1','1','1','1','1','1','0','0','1','1','1','1','1','0','0','0','0','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','1','1','1','1','1','0','0','0','0','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','0','0','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','0','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','1','1','0','0','1','1','1'),
('0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0'),
('0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));

constant PokemonString : PokemonBits := 
(("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000101","010101","010101","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","000101","000001","000101","010110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000101","000001","010110","010110","000110","010110","000101","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","000101","000101","010110","010110","010110","000110","010110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010101","000001","000101","000110","000110","010110","000110","000110","010110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000001","010110","010110","000110","010110","010110","000110","000101","010110","000110","000101","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000101","000110","000110","000110","010110","010110","010101","011010","010101","000101","010110","010110","000101","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000101","000110","010110","010110","010110","010110","010101","011001","101001","011001","010101","010101","010110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011011","000110","000110","010110","000110","010110","010110","010101","101001","101001","101001","101001","010101","010101","010110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000110","000110","000110","000110","000110","010110","010101","100101","111001","111001","101000","101000","101001","010101","010110","010110","010110","000110","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000110","000110","010110","000110","000110","010110","010101","010101","101001","111101","111100","111000","111000","101000","101001","010101","010110","000110","010110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","000110","000110","000110","000110","000110","000110","010110","010101","111001","111101","111100","111100","111000","111000","101000","101001","010101","010101","010110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","000101","000110","000110","000110","010110","010101","010101","101001","111100","111100","111100","111100","111100","111000","101000","101001","101001","010110","010110","000110","010110","010110","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","011010","000110","000110","000110","000110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111000","111000","101000","101001","010110","010110","010110","010110","010110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000110","000110","000110","000110","010110","010101","010101","101001","111101","111100","111100","111100","111100","111100","111101","111101","111101","101001","010101","010101","010110","010110","010110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000000","000000","000000","000000","101010","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000110","000110","000110","000110","000110","010110","010101","100100","111001","111100","111100","111100","111100","111100","111101","111001","101001","010101","010101","010101","000101","000110","010110","010110","010110","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","010110","010101","010101","000000","000000","101011","010101","010101","000101","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000110","000110","000110","000110","000110","010110","010101","010101","111101","111101","111000","111100","111100","111101","111001","101001","010101","010101","010101","010110","000110","000110","000110","010110","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","010110","000101","010110","010110","010110","000110","000000","010110","000101","000101","000001","010110","010110","000101","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011011","000110","000110","000110","000110","000110","000110","010101","010101","111001","111101","111000","111101","111101","111001","101001","010101","010101","010101","000101","000101","010110","000110","000110","011010","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","011010","010110","000101","000110","010110","010110","010110","000110","000110","010110","010110","000001","000010","000110","000110","010110","000110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011011","000110","000110","000110","000110","000110","010110","010110","010101","101001","111101","111101","111101","111101","101001","010101","010101","010101","010101","010110","010110","010110","000110","011010","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010101","010101","000101","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010101","010101","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","101011","011010","010110","010110","010110","010110","010110","010110","010110","010110","010110","101010","101011","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","011010","010110","010110","000110","000110","010110","000110","000110","000110","000110","000110","000110","010110","000110","010110","000110","000110","010110","000110","000110","010110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000110","000110","000110","000110","000110","010111","000110","010101","101010","111110","111101","101001","101001","010101","010101","010110","010110","010110","010110","010110","010110","011010","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","000001","000101","010110","010110","010110","010110","010110","010110","000110","010110","010110","010110","010110","010110","010110","010110","010110","010110","000101","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","101010","011010","010110","010110","010110","010110","010110","000110","000110","010110","010110","010110","000110","000110","010110","010110","010110","010110","010110","000110","000101","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","010110","010110","010110","010110","000110","010110","010110","000110","000110","000110","010110","010110","000110","000110","000110","000110","000110","000110","010110","000110","000110","010110","000110","010110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","000110","000110","000110","000110","000110","000110","010110","000101","011001","101010","101001","010101","010101","000101","010110","010110","010110","010110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","101011","101011","101011","101011","101010","101010","101011","101010","101010","101010","101011","101011","101011","011010","010110","000101","000101","000110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010110","010110","010110","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","010110","010110","010110","010110","010110","010110","000110","000110","000110","010110","010110","010110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010110","000110","010110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","010110","010110","000110","010110","010110","010110","000110","000110","000110","000110","000110","010110","000110","000110","000110","000110","010110","000110","000110","000010","000110","010110","000110","000110","000110","010110","010110","010110","010110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","000101","000110","000110","000110","000110","000110","000110","010110","010110","000101","010101","010101","000101","000101","000110","000110","000110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","011010","010110","000101","000110","010110","010110","010110","010110","010110","010110","010110","010110","000110","000110","000110","010110","000110","010110","000110","010110","000110","000110","000110","000110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","010110","010110","010110","010110","000110","000110","010110","010110","010110","010110","000110","000110","000110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","000110","010110","010110","010110","010110","010110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","101011","010110","010101","010101","010110","010110","000110","010110","010110","010110","010110","000110","010110","010110","010101","010101","010101","010110","010110","000110","000110","000110","000110","000110","000110","010110","000110","010110","010110","010101","010101","010110","010110","010110","010110","000110","011010","000000","000000","000000","000000","000000","000000","000000","000000","010110","000001","000101","000001","000001","000101","000110","000110","010110","000110","000110","010110","010110","010110","010110","000110","000110","000110","000110","011011","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000001","000001","000110","010110","010110","000110","000110","000110","000110","010110","010110","010110","010110","010110","010110","010110","000110","010110","010110","000110","000110","000110","000110","010110","010110","010101","010101","010101","010101","010101","010101","010101","010101","010101","010110","010110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","010110","010110","010110","010110","010110","000110","000110","010110","010110","010110","010110","010110","010110","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010110","010110","000110","010110","010110","010110","010110","000110","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","010101","010110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010101","010101","010101","010101","010101","101001","101001","010110","010110","010110","000110","010110","000110","000110","000110","000110","000110","010110","010101","010101","101001","010101","010101","010110","010110","010110","000101","011010","000000","000000","000000","000000","000000","000000","101010","000101","000001","000001","000001","000001","000110","000110","000110","000110","000110","010110","010110","010110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","011010","101011","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000001","000001","000010","010110","010110","010110","000110","010110","000110","000110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","000110","000110","000110","000110","010110","010110","010101","101001","101001","101001","101001","101000","101000","101001","101001","010101","010110","010110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","000001","010110","010110","010110","101010","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","010110","010110","010110","010110","000110","000110","010110","010110","010110","010110","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","101001","101001","101001","101001","101001","101001","101001","101001","010101","010101","010101","010101","010101","010101","010110","000110","010110","000110","000110","010110","010110","000110","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","000101","000101","010110","000110","000110","010110","010110","010110","010110","010110","010110","010101","010101","010101","010101","011001","101001","101001","101001","101001","101001","101001","010101","010110","010110","010110","000110","000110","000110","000110","000110","010101","010101","101001","101001","101001","010101","010101","010110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","101010","000001","000001","000001","000001","000001","000110","000110","000110","010110","010110","010110","010110","010110","000110","000110","000110","000110","010110","010110","010110","000110","000110","000110","000110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000101","000001","000010","000010","010110","010110","010110","000110","010110","010101","010101","010101","010101","010101","010101","010101","010110","010101","010101","010101","010101","000110","000110","000110","000110","010110","010101","101001","111000","111000","111000","111000","111000","111000","101000","101000","010101","010101","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","000001","000001","000001","010110","000110","010110","010110","010110","010110","010110","011010","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","010110","000110","010110","000110","000110","000110","000110","000110","000110","000101","010101","010101","010101","010101","100101","101001","101001","101001","101001","101001","101001","101000","101000","101000","101000","101000","101000","101000","101000","101000","101001","101001","101001","101001","101001","010101","010101","010101","010101","010110","010110","000110","000110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","000101","000001","000001","010110","000110","010110","010110","010110","010110","010110","010101","010101","010101","010101","100100","101000","101000","101000","111000","111000","111100","111000","101001","101001","010101","010110","010110","010110","000110","000110","000110","010110","000101","010101","101001","101000","101000","101001","101001","010101","010101","010110","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","010110","000001","000001","000001","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","000110","000110","000110","010110","010110","010110","010110","010110","010110","010110","000110","010110","101010","000000","000000","000000","000000","101111","000101","000101","000110","000110","000110","010110","010110","010110","010101","101001","101001","101001","101001","101000","101001","101001","101001","101001","101001","101001","101001","010110","000110","000110","000110","010110","010101","111001","111100","111100","111100","111100","111100","111000","111000","101000","010101","010101","000110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010101","000001","000001","000001","000110","000110","010110","010110","000110","000110","000110","010110","010110","010110","000101","010110","011010","101010","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000110","010110","010110","010110","000110","010110","010110","010110","010101","010101","010101","010101","010101","101001","101001","101001","101000","101000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","101000","101000","101001","101001","010101","010101","010101","010110","010110","010110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","000001","000101","000101","000001","000001","010110","010110","010110","010110","010110","010101","100101","101001","101001","111001","111000","111000","111100","111100","111100","111100","111100","111000","111000","101001","010101","010110","010110","010110","000110","010110","000110","000110","010101","101001","111101","111000","111000","101000","111001","101001","010101","010101","010110","010110","010110","010110","000110","101011","000000","000000","000000","000000","000000","010110","010110","000110","010110","010110","010110","000110","000110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010101","010101","010101","010101","010101","010110","010110","000110","010110","000110","000101","010110","101011","000000","000000","101011","000101","000101","000110","000110","000110","010110","010110","010101","010101","101001","101001","101000","101000","101000","111000","101000","101000","101000","101000","101000","101001","010101","000101","010110","010110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","000110","010110","010110","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000001","000101","000101","000001","000010","010110","000110","000110","000110","010110","010110","010110","010110","000110","010110","000110","000110","000110","000110","010110","010110","011010","101011","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","010110","010110","000110","000110","000110","000110","010110","010110","010101","000101","010101","010101","101001","101001","101001","111001","111000","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","111000","111000","111000","111000","101000","101001","100101","010101","010101","010101","010110","010110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","000101","000001","000001","000101","000110","010110","010110","010110","010101","101001","101001","101001","111001","111000","111000","111000","111000","111100","111100","111100","111100","111100","111000","111000","101001","010101","010110","010110","010110","010110","010110","010110","010101","101001","111101","111101","111100","111000","111000","111000","101000","101001","010101","010101","010110","000110","010110","000110","010110","101011","000000","000000","000000","000000","010110","010110","010110","010110","010110","010110","010110","010110","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010110","010110","010110","000110","010110","010110","000110","000101","101010","000000","011010","000001","000101","000101","000110","000110","010110","010110","010101","010101","111001","111100","111000","111100","111000","111000","111000","111000","111100","111000","111000","101001","010101","010101","010110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","000110","010110","010110","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000101","000001","000001","000010","010110","000110","000110","010110","010110","010110","010110","010110","010110","010110","010110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","101010","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","000110","010110","000110","010110","000110","000101","010101","010101","010101","010101","101001","101001","101000","111000","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","101000","101000","101001","101001","010101","010101","010110","010110","000110","010110","000110","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","000001","000101","000101","000110","000110","010110","010110","010110","010101","101001","111101","111001","111101","111100","111000","111000","111000","111100","111100","111100","111100","111100","111000","111000","101001","010101","010110","010110","000110","010110","010110","010101","010101","111001","111101","111100","111100","111100","111000","111000","101000","101000","101001","010101","010101","010110","010110","000110","010110","010110","101011","000000","101010","010110","010110","010110","010110","010110","010110","010101","010101","010101","010101","010101","100101","101001","101001","101001","101001","101001","101001","101001","101001","101001","101001","100101","010101","010101","010101","000101","010110","000110","010110","010110","010110","010110","010110","000001","000101","000101","000110","000110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010110","010110","010101","100101","111101","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000001","000001","000001","000010","000110","000110","000110","000110","000110","010110","010101","010101","010101","010101","010101","010101","010101","000110","010110","010110","010110","010110","000110","000110","010110","010110","010110","010110","010110","010101","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","101111","011010","000110","000110","010110","000110","010110","000110","010110","010101","010101","010101","101001","101001","101000","111100","111100","111000","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","101000","111001","101001","010101","010101","010110","010110","000110","010110","000110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","000101","000110","000110","000110","000110","010110","000110","000110","010101","101010","111110","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101001","010101","000101","000110","000110","010110","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111000","101000","111001","101001","010101","010110","010110","010110","000110","000110","010110","000110","000110","010110","000110","000110","000110","010110","010101","010101","010101","011000","101000","101000","101000","111000","111000","111000","111000","111000","101000","101000","101000","111001","111001","101001","101001","101001","011001","010101","000101","010110","010110","000110","000110","010110","010110","000010","000101","000101","000110","000110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101001","010101","010101","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000101","000110","000001","000110","010110","000110","000110","010101","101001","101001","101001","100101","010101","010101","010101","010101","010101","010101","010101","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","101011","000000","000000","101010","101010","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","101010","010110","000110","000110","010110","000110","010110","010110","010101","010101","010101","101001","101001","111000","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101000","101001","010101","010101","000110","000110","010110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000101","000001","000110","000110","010110","000110","000110","010101","101010","101010","101001","101000","100100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101001","010101","000101","000110","000110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","101001","010101","010101","010110","010110","010110","010110","000110","010110","000110","000110","010110","010110","010101","010101","101001","101001","111000","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","101000","101000","101000","101001","101001","010101","010101","010101","010110","010110","010110","010110","000110","000110","000101","000110","000110","000110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101001","010101","010101","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000001","000101","000001","000110","000110","000110","000110","010101","101001","101001","101000","101000","101000","101001","101001","101001","101001","010101","010101","010101","010101","010101","010101","010101","010101","010110","010110","000110","000110","011010","101011","010101","000101","010110","010110","010110","010101","010110","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","010110","000101","000110","000110","000110","000110","010110","010101","010101","010101","101001","111001","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101000","101001","011001","010101","010110","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000101","000110","000110","000110","000110","000110","000110","010110","010110","010101","010101","010101","010100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101001","010101","000101","000110","010110","010101","101001","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","101000","101001","010101","010101","010101","010110","000110","000110","010110","010110","000110","010101","010101","101001","101001","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","101000","101000","101001","101001","010101","010101","010110","010110","010110","010110","000110","000110","000110","000110","010110","010110","010101","111110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","101001","010100","010101","010101","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","010101","010101","010110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000101","000001","000110","000110","010110","000110","000101","010101","101001","111001","111000","111000","101000","101000","101000","101000","101000","101000","101001","101001","101001","101001","010101","010101","010101","010101","010110","010110","000110","000110","000101","000001","000101","010110","010110","010110","010110","010110","010110","010110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","101011","000101","010110","000110","000110","000110","010110","000110","010101","010101","101001","111001","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","101001","010101","010101","010110","000110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010101","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","000101","010110","010101","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","101000","101001","010101","010101","010110","000110","000110","010110","010110","000101","010101","101001","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111100","111100","111100","111100","111100","111100","111100","111000","101000","101000","101001","101001","010101","000101","010110","010110","010110","000110","000110","000110","000110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","101000","010100","010101","010101","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000110","000101","000101","000110","000110","000110","010110","010101","101010","111101","111101","111100","111100","111000","111000","111000","111000","111000","101000","101000","101000","101000","101001","101001","101001","010101","010110","000110","000110","000110","000101","000101","000110","010110","010110","010110","010110","000110","000110","000110","000110","010110","010110","010110","010110","010110","101010","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","101011","000001","000101","000110","010110","000110","000110","010110","010110","010101","101001","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","101000","101001","010101","010101","010110","010110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010101","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010101","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","101001","011001","010110","000110","010110","010110","010110","010101","010101","101001","111101","111100","111100","111100","111100","111000","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","101000","101001","011001","010101","010110","010110","010110","000110","000110","000110","000110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","101000","101001","010101","010101","100100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000101","000110","000101","000110","010110","000110","000110","000101","010101","101001","101001","111001","111101","111100","111100","111100","111100","111100","111000","111000","111000","111000","101000","101001","101001","010101","010110","000110","000110","000110","000110","000110","000110","010110","010110","000110","010110","010110","010110","000110","000110","000110","010110","010110","010110","010110","010110","010110","010110","010110","101010","101111","000000","000000","000000","000000","000000"),
("000000","101011","000000","000101","000001","000110","000110","000110","010110","010110","010101","101010","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","101000","101001","010101","010110","010110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010110","010110","010110","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","101000","101001","010101","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111001","101001","010101","000110","000110","010110","010110","010101","010101","111001","111100","111100","111100","111100","111000","111100","111100","111101","111101","111101","111101","101001","101001","101001","111101","111101","111100","111100","111100","111100","111100","111100","111000","111100","111100","111000","101000","101001","101001","010101","000110","010110","010110","000110","000110","000110","000110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101001","010101","010101","010110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000101","000110","000101","000110","000110","000110","010110","000110","010101","010101","010100","101000","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010110","010110","000110","000110","000110","000110","000110","010110","000110","010110","010110","010101","010101","010101","010101","010110","010110","010110","010110","010110","010110","010110","010110","000110","000110","010110","010110","011010","101010","000000","000000"),
("101011","000001","000001","000001","000001","000110","010110","010110","010110","000110","010101","101001","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","101001","010101","010101","010110","010110","010110","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010110","010110","010110","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","101000","101001","100101","010100","010100","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","010101","000110","010110","010110","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111101","111001","101001","010101","010101","010101","010101","010101","010101","010101","101001","111101","111101","111100","111100","111100","111100","111100","111000","111000","111001","101001","010101","010101","010110","000110","000110","000110","000110","000110","000110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101001","010101","010101","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000101","000110","000110","000110","000110","000110","010110","010110","010110","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","101001","010101","010101","010110","000110","000110","000110","000110","000110","000110","010101","010101","101001","101001","101001","010100","010100","010100","010101","010101","010110","010110","010110","010110","000110","000110","000110","000110","000101","010101","101010","000000","000000"),
("000101","000001","000001","000001","000001","000001","000110","000110","010110","010110","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101000","101001","010101","010110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111000","111001","100100","010100","111001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","010101","000110","000110","000110","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111101","101001","100101","010101","010101","010101","010110","010110","010110","010110","010101","010101","101001","101000","111100","111100","111100","111100","111100","111100","111101","111001","010101","010101","010110","000110","010110","000110","000110","000110","000110","000110","010110","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010101","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000101","000110","000110","000110","000110","000110","000110","000110","000110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","000110","000110","000110","000110","000110","000110","010110","010101","010101","101001","101000","101000","101000","101001","101001","101001","100101","010101","010101","010101","010101","010110","010110","010110","010110","010110","010101","101111","000000","000000"),
("101111","000101","000001","000001","000001","000001","000101","000110","000110","010110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","101001","010101","010110","000110","010110","000101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000101","000101","000110","000110","000110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","100100","101000","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111001","100101","010101","010110","000110","000110","000110","010101","100101","111001","111101","111100","111100","111100","111100","111100","111101","101001","010101","010101","010110","010110","010110","010110","010110","010110","010110","010110","010101","010100","101000","111100","111100","111100","111100","111100","111101","111001","101001","010101","010110","010110","000110","010110","000110","000110","000110","000110","010110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","101001","010101","010101","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","000110","000110","000110","000010","000110","000110","000110","000110","000110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010110","010110","000110","000110","000110","010110","010101","010101","101001","111001","111000","111000","111000","111000","111000","101000","101000","101001","101001","101001","011001","010101","000110","000110","010110","010110","010110","000000","000000","000000"),
("000000","010110","000001","000001","000001","000001","000001","000110","000110","000110","010110","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","111101","111001","101001","101000","111001","111101","111101","111100","111100","111100","111100","111100","111100","111000","111000","111100","111100","111000","101000","101001","010101","010110","010110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010101","000101","000110","000110","000110","000110","000001","000001","000001","000110","000110","010110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","111100","111100","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111001","010101","010101","010110","000110","000110","000110","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","101001","010101","010101","010110","010110","010110","010110","011010","011010","010110","010110","010110","010101","010101","101001","111100","111100","111100","111100","111101","111001","100101","010101","010110","010110","000110","010110","000110","000110","000110","000110","000110","010110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","100100","100100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","101000","010101","010101","010110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","101011","011010","010110","010110","010110","010110","000101","000110","000110","000110","000110","000010","000001","000001","000110","000110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010100","010101","000110","000110","000110","000110","010110","010101","010101","101001","111101","111100","111100","111000","111000","111000","111000","111000","101000","101000","101001","101001","010110","010110","010110","010110","010110","101010","000000","000000","000000"),
("000000","000000","000101","000001","000001","000001","000001","000110","000110","000110","000110","010110","010101","010101","111001","111101","111100","111100","111100","111100","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","101001","011001","010101","010101","010101","010101","010101","010101","011001","101001","111101","111101","111100","111100","111100","111100","111000","111000","111100","111000","101000","101001","010101","010110","010110","010110","000110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","101011","101111","000000","101111","000001","000001","000001","000001","000110","000110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111101","010100","010101","010110","010110","000110","000110","000110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111001","101001","010101","010110","010110","101010","101111","000000","101111","101011","010110","000110","010110","010101","101001","111101","111100","111100","111100","111101","111101","100101","010101","010101","010110","010110","010110","010110","000110","000010","000110","000110","000110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","100100","101000","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","000110","000110","010110","101010","000000","000000","000000","000000","101011","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","000110","000110","000110","010110","000110","000110","000110","000110","010110","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101000","010101","010101","000110","000110","000110","000110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111001","101001","010101","010110","010110","010110","010110","000000","000000","000000","000000"),
("000000","000000","101010","000001","000101","000001","000001","000110","000110","000110","000110","010110","010110","010101","101001","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","010101","010101","010110","010110","010110","000110","010110","010110","010101","010101","101001","111101","111101","111100","111100","111100","111000","111000","111100","111100","101000","101001","010101","010110","010110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","000001","000001","000001","000001","000110","000110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111000","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010101","010101","010110","000110","000110","000110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111000","101001","010101","010101","000110","101011","000000","000000","000000","000000","101011","000110","010110","010101","101001","111101","111100","111100","111100","111100","111101","100101","010101","010110","010110","010110","000110","010110","010110","000010","000001","000110","000110","000110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010110","010110","000110","011010","000000","000000","101010","010110","000110","000110","010110","010110","010110","000110","010110","010110","000110","000110","000110","010110","010110","010110","010110","000110","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","010101","010101","000110","000110","000110","000110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","100101","010101","010110","010110","010110","010110","000000","000000","000000","000000"),
("000000","000000","000000","010101","000001","000101","000001","000101","000101","000110","000110","000110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010110","000110","000110","010110","010110","000110","000110","010110","010101","010101","100101","111101","111100","111100","111100","111100","111100","111100","111100","101000","101001","010101","010110","000110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","101011","101011","101010","101010","101010","101010","101011","000110","000110","000010","000001","000110","000110","010110","010110","010101","100101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010100","010101","010101","010110","010110","000110","010110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111000","101001","010101","000101","010110","000000","000000","000000","000000","101111","000101","010110","010101","101001","111001","111100","111100","111100","111100","111001","101001","010101","010110","000110","000110","000110","010110","000110","000001","000001","000001","000110","000110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010110","000110","000110","010110","101011","010110","000101","010110","010110","000110","000110","010110","010110","010110","010101","010101","010101","010101","010110","010110","010110","010110","000110","010110","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","000110","000110","000110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010101","010101","010110","010110","000110","101011","000000","000000","000000","000000"),
("000000","000000","000000","101111","000001","000101","000001","000101","000101","000110","000110","000110","010110","010110","010101","100101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101001","010101","010110","000110","000110","010110","010110","010110","010110","010110","010110","010101","010101","101001","111100","111100","111100","111100","111100","111100","111100","101000","101001","010101","010110","010110","000110","010110","101011","000000","000000","000000","000000","000000","011010","010110","010110","000110","010110","000110","010101","000101","000101","010110","000110","000110","000110","000110","000110","000110","000110","010110","010101","100100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","101001","010101","010110","000110","010110","000110","010110","010110","010110","010110","010101","111001","111100","111100","111100","111100","111100","111100","101000","101001","010101","010110","011010","000000","000000","000000","101011","010101","010101","010101","011001","111101","111100","111100","111100","111100","111101","101001","010101","010110","010110","000110","000110","000110","010110","000110","000001","000001","000001","000110","000110","010110","010110","010101","111001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101001","010101","000110","000110","000110","000110","000110","000110","010110","000101","010101","010110","010110","010101","010101","010101","010101","010101","011001","101001","100101","010101","010101","010101","010101","010110","010110","010110","000110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010110","000110","000110","010110","010101","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010101","010110","010110","010110","101111","000000","000000","000000","000000"),
("000000","000000","000000","000000","010110","000001","000010","000010","000101","000101","000110","000110","010110","010110","010110","010101","101001","111101","111100","111100","111100","111101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010110","000110","000110","011010","011010","011010","010110","010110","010110","010110","010110","100100","111101","111100","111100","111100","111100","111100","111100","111000","101001","010101","010110","010110","000110","010110","000000","000000","000000","101011","010110","000101","000110","010110","000110","000110","000110","010110","010110","010110","000110","010110","000110","000110","000110","000110","000110","000110","000110","000101","010101","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010101","010110","010110","010110","000110","010110","010110","000110","010110","010110","010101","111101","111100","111100","111100","111100","111100","111100","101000","011001","010101","010110","011011","000000","000000","000000","010110","000101","010101","010101","111101","111100","111100","111100","111100","111001","101001","010101","010101","010110","010110","000110","000110","000110","000110","000110","000110","000010","000010","000110","000110","000110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","010101","010110","010110","000110","000110","000110","010110","010110","010101","010101","010101","010101","101001","101001","101001","101000","101000","101000","101000","101000","101001","101001","101001","011001","010101","010101","010110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010101","010110","000110","010110","010101","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010101","010110","010110","010110","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000101","000110","000110","000101","000101","000110","000110","000110","010110","010110","010101","010101","101001","111101","111101","111000","111001","101001","101000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","010101","010101","000110","000110","101111","101111","101010","010110","011010","010110","010110","010101","010100","111101","111100","111100","111100","111100","111100","111100","101000","101001","010101","000101","010110","000110","000110","101111","101011","010110","010110","010110","010110","010110","010101","010101","010110","010110","010101","010101","010101","010101","010101","010110","000110","000110","000110","010110","010110","000110","000110","010101","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111001","101001","010101","010110","010110","000110","000110","011010","101111","000110","000110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","101000","011001","010101","010110","011010","000000","000000","010110","010110","010101","010101","111101","111101","111100","111100","111101","111101","101001","010101","010101","010110","010110","000110","000110","000110","000110","000110","010110","010110","000110","000110","000110","000110","000110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","010101","010110","010110","000110","000110","010110","010101","010101","010101","100101","101001","101001","101001","101001","111000","111100","111000","111000","111000","111000","111000","111000","101000","101000","101001","010101","010101","010101","010110","010101","010101","101000","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101000","010101","010101","010110","010110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","010101","010101","010110","010110","010110","101010","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","101010","000110","000110","000110","000101","000101","000110","000110","000110","010110","010110","010101","101001","111110","111101","101001","100101","010101","010100","101000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101001","010101","000110","000110","101010","000000","000000","101010","010110","010110","010110","010101","010101","101001","111100","111100","111100","111100","111100","111100","101001","100101","010101","010110","000110","010110","000110","011011","000110","010110","000110","000110","010110","010110","010101","010101","010101","010101","010101","010101","101001","011001","010101","010101","010101","010101","010101","010110","010110","010110","010110","010101","010101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111001","101001","010101","010110","010110","010110","010110","011010","000000","101111","000110","000110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","101000","101001","010101","010110","010110","000000","011010","000101","010101","010101","101001","111101","111100","111100","111100","111101","101001","010101","010101","010110","010110","010110","010110","010101","010101","010101","010110","010110","000110","010110","000110","000110","000110","000110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111100","111000","101001","010101","010101","000110","000110","010110","000101","010101","010101","101001","101001","111101","111101","111110","111001","101001","101000","101000","111000","111100","111000","111000","111000","111000","111000","101001","101001","010101","010101","010110","010110","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","010101","010101","010110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010101","010110","010110","010110","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000101","000110","000110","000101","000101","000110","000110","000110","000110","000110","010110","010101","101001","010101","010101","010101","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101001","010101","010110","010110","010110","000000","000000","000000","011010","010101","010110","010110","010101","101001","111100","111100","111100","111100","111100","111100","101001","010101","010101","010110","000110","000110","000110","000110","000110","000110","010110","010110","010101","010101","100101","101001","101001","101001","101001","101000","101000","101000","101000","101001","101001","101001","010101","010101","010101","010110","010110","010101","010101","111010","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","101001","010101","010101","010110","000110","010110","011010","000000","000000","101111","000110","000110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111000","101001","010101","010101","010110","010110","010110","010101","010101","101001","111101","111100","111100","111100","111101","101001","010100","010101","010110","010110","010110","010101","010101","101001","011001","010101","010101","010110","010110","010110","000110","000110","000110","000110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","101001","010101","010110","010110","000110","010101","010101","101001","101001","111101","111101","111101","101001","101001","010100","010100","101000","101000","111000","111100","111100","111100","111000","111000","111000","101000","111000","101001","010101","010101","010110","010110","010101","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","101111","000101","000101","000110","000101","000110","000110","000110","000110","000110","010110","010110","010101","010101","010110","010110","010110","010101","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","101001","010101","010101","010110","010110","000000","000000","000000","010101","010110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111000","101001","010101","000101","010110","000110","000110","010110","000110","010110","010101","010101","010101","101001","101001","111000","111000","111000","111000","111000","111000","111000","101000","101000","111000","101000","101000","101001","101001","010101","010101","000101","010110","010101","010101","111001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","010101","010110","010110","000110","011010","000000","000000","000000","000000","000110","010110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111000","101000","011001","010101","010110","010110","010101","010101","101001","111101","111100","111100","111100","111101","101001","010100","010101","010101","010110","010101","010101","100101","101001","101001","101001","100101","010101","010101","010110","010110","010110","000110","000110","000110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111001","010100","010101","010110","010101","010101","010101","101001","111101","111101","111101","111101","101001","010101","010101","010100","101001","101000","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101000","101001","010101","010101","010110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010110","010110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","010101","010110","010110","000110","000110","101011","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010110","000110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010110","010110","101011","000000","000000","011010","010101","010110","010110","010101","111001","111100","111100","111100","111100","111100","111001","100101","010101","010110","000110","000110","010110","010110","010110","010101","010101","011001","101001","111001","111000","111100","111101","111101","111101","111101","111100","111100","111100","111100","111000","111000","101000","111000","101000","101001","010101","010101","010101","010101","010101","101001","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","010101","010101","010110","000110","010110","000110","010110","101011","101111","000000","000000","010110","010110","010110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111000","111000","101000","010101","010101","010101","010101","101001","111101","111100","111100","111100","111101","101001","010101","010100","010101","010101","010101","010101","101001","111001","101000","101000","101000","101001","100101","010101","010101","010110","000110","000110","000110","000110","010110","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111001","101001","010101","010110","010110","010101","010101","101001","111101","111101","111101","111101","101001","010101","010110","010101","101001","101000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101000","101001","010101","010110","010110","010101","100101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010101","010110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","010101","010110","000110","010110","010110","101111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","101111","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","000110","010110","010110","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","101001","010101","010110","010110","010110","000000","000000","011010","000110","010110","010101","010101","111101","111100","111100","111100","111100","111101","101001","010101","010101","000110","000110","010110","010110","010101","010101","100101","101001","111001","111100","111101","111101","111101","111001","101001","100100","100100","101000","111000","111100","111100","111100","111100","111000","111000","101000","111001","101001","010101","010101","010101","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","010100","010100","010101","010110","010110","000110","010110","010110","010110","000101","010110","101011","010110","010110","000110","010110","010101","111001","111100","111100","111100","111100","111100","111100","111100","111000","101000","100101","010101","010100","101001","111101","111100","111100","111100","111100","101001","010100","010101","010101","010101","010100","100100","101001","111101","111100","111100","111000","111000","111000","101001","101001","010101","010101","000101","000110","010110","000110","010101","100101","111001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101000","010101","010101","010110","010101","010101","101001","111101","111101","111100","111101","101001","010101","010110","000110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111000","111100","111100","111000","101000","101000","101001","010110","010110","010101","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101000","010101","010101","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","100101","010101","010110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","011010","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010110","010110","010110","000000","101111","011010","010110","010110","010101","101001","111101","111100","111100","111100","111100","111001","100101","010101","010110","000110","000110","010110","010110","010101","100101","111001","111101","111101","111100","111100","111001","101001","010101","010101","101001","101000","111000","111100","111100","111100","111100","111100","111100","111100","101000","111000","101001","101001","010101","010101","010110","010101","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","010100","010101","010101","010101","010110","010110","000110","010110","010110","010110","010110","000110","000110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111000","111000","111000","101000","101000","111101","111100","111100","111100","111100","111000","100100","010100","010101","100101","100101","101000","111001","111100","111100","111100","111100","111100","111000","111000","111000","101000","101001","010101","010101","000110","000110","000110","010110","010101","100101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","011001","000101","010101","010110","010101","101001","111101","111100","111100","111100","111000","010101","010101","010110","000110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","101000","101000","111100","111100","111100","111000","101000","101001","010101","010110","010101","010101","101000","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010101","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010101","010110","010110","010110","010110","101010","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","010101","010101","010110","010110","101011","011011","010110","010110","010110","010101","111001","111100","111100","111100","111100","111101","101001","010101","010101","000110","000110","000110","010101","010101","101001","111001","111100","111100","111100","111101","101001","100101","010101","010101","100101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","101001","101001","010101","010101","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101000","101000","101001","010101","010101","010101","010101","010110","010110","010110","010110","010110","010110","000110","000110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111000","111000","111000","111000","111100","111100","111100","111100","111100","111000","111000","101000","101000","101000","101000","111001","111101","111100","111100","111100","111100","111100","111100","111100","111000","101000","101000","111001","101000","010101","010101","000110","000110","010110","010110","010101","100101","111000","111100","111100","111100","111100","111100","111100","111100","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","010101","010101","010110","010101","010101","111001","111101","111100","111100","111000","101000","010101","010110","000110","000110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111000","101000","100100","111000","111100","111100","111000","111000","101000","010101","010101","010101","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010101","010100","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010101","010110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000101","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","101001","010101","010110","010110","010110","010110","000110","010101","010101","101001","111101","111100","111100","111100","111100","111001","010101","010101","000110","000110","010110","000110","010101","101001","111101","111101","111100","111100","111100","101001","101001","010101","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111000","111100","111000","111000","101000","101001","010101","010101","010101","010101","010101","111101","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","111000","111000","101001","101001","101001","010101","010101","010101","010101","010110","010110","000110","000110","000110","000110","010101","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","101001","101001","010110","000110","000110","010110","010110","010101","010100","101000","111100","111100","111100","111100","111100","111100","111000","101000","111000","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111001","010101","010101","010110","010101","010101","101001","111101","111100","111100","111100","111000","101000","010101","010110","000110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","101000","101000","010100","111000","111100","111100","111000","111000","101000","010101","010101","010101","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010101","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","100101","010101","010110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000101","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010101","011001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010110","010110","000110","000110","000110","010101","101001","111001","111100","111100","111100","111100","111101","101001","010101","010110","000110","010110","000110","010101","100101","111001","111101","111100","111100","111100","111101","011001","010101","010110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","111101","111100","111000","111000","101000","101001","010101","010101","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","111000","101000","101000","101001","101001","101001","010101","010101","010101","000110","000110","000110","000110","000110","010101","100101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","011001","010110","000110","000110","000110","010110","010101","100100","111000","111100","111100","111100","111100","111100","111000","111000","100100","101000","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010101","010110","010101","010101","111001","111100","111100","111100","111100","111000","101000","010101","000110","000110","010110","010110","010101","011001","101001","111101","111101","111101","111101","111001","101001","010101","010100","101000","111100","111100","111000","111000","101000","101001","010101","010110","010101","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101001","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","010101","010110","000110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","000101","000110","000110","000110","000101","000101","000101","000110","000110","000110","000110","000110","000110","000110","000110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010101","010110","010110","000110","010101","010101","111101","111100","111100","111100","111100","111101","111001","010101","010101","010110","010110","010110","010101","010101","111001","111101","111000","111100","111100","111100","101000","010101","000101","000110","000110","010101","101001","111100","111100","111100","111100","111100","111100","111100","101000","101000","100100","111001","111100","111100","111000","101000","101001","010101","010101","010101","010101","010101","111101","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","101000","101000","101000","101001","101001","010101","010101","010101","000101","000110","000110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111100","111100","111100","111100","111100","111100","111100","111101","111001","010101","010101","010110","010110","010110","010101","010101","010101","111101","111100","111100","111100","111100","111100","111100","111000","101001","010100","010100","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","100101","010101","010110","010101","010101","101001","111101","111100","111100","111100","111000","111000","101001","010101","010110","010110","000110","010110","010110","000101","010101","101001","101001","101001","101001","100101","010101","010101","010101","111001","111100","111100","111100","111000","101000","101001","010101","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","010101","010100","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","010101","010110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","000101","000101","000101","000101","101011","010110","000101","000110","000101","000110","000110","000110","000110","000110","010110","010101","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101001","010101","010101","000101","010101","101001","111001","111100","111100","111100","111100","111101","111001","100101","010101","010101","010110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111000","101001","010101","010110","000110","000110","010101","101001","111001","111101","111100","111100","111100","111100","111100","101000","101001","010100","101001","111101","111100","111000","111000","101001","100101","010101","000110","000101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","111000","101000","101000","101000","101001","011001","010101","000101","010110","010110","010101","010101","111001","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111001","100101","010101","010110","000110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","101000","101001","010100","010100","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","101000","111100","111100","111100","111100","101001","010101","010101","010110","010101","010101","111101","111100","111100","111100","111100","111000","111000","101000","010101","010101","010110","010110","000110","000110","000110","000110","010101","010101","010101","010101","010101","010101","010101","010101","111101","111100","111100","111100","111000","101000","101001","010101","010110","010110","010101","101001","111100","111000","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","100100","010100","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","010101","010110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010101","010110","000000","000000","000000","101111","000101","000110","000001","000101","000110","000110","000110","000110","010110","010101","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","010100","010101","010101","101001","111101","111101","111100","111100","111100","111101","111001","100101","010101","010101","010110","000110","010110","010101","010101","111001","111100","111100","111100","111100","111100","101000","101001","010101","010110","000110","000110","000110","010101","101001","111101","111101","111100","111100","111101","111101","101001","010101","010100","101001","111101","111100","111100","111000","101000","101001","010101","000110","000101","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","111000","101000","101000","101001","011001","010101","010101","010110","010110","010101","010101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","101001","010101","010101","010110","010110","000110","010110","010110","101001","111001","111101","111100","111100","111100","111100","111100","111100","111100","101000","101001","010101","010101","010101","111001","111100","111100","111100","111100","111100","111100","111100","101000","010100","111100","111100","111100","111000","101001","010101","010101","010110","010101","010101","111101","111100","111100","111100","111100","111000","111000","101000","101001","010101","010101","010110","010110","000110","000110","000110","000110","000110","000110","010110","010110","010101","010101","101001","111101","111100","111100","111100","111000","101000","101001","010101","010110","010110","010101","101001","111101","111100","111100","111000","111000","111100","111100","111100","111100","111100","111000","101000","101000","100100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","010101","010101","010110","000110","000110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000101","000101","000110","000110","000110","000110","000110","010110","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","100100","101000","101001","111101","111100","111100","111100","111100","111101","111001","101001","010101","010101","010110","000110","000110","010110","010101","101001","111101","111100","111100","111100","111100","111100","101000","101001","010101","010110","000110","000110","000110","010110","010101","101001","101001","111101","111101","101001","101001","010101","010101","010100","101001","111100","111100","111100","111000","101000","101001","010101","000110","010110","010101","111001","111100","111100","111100","111100","111100","111100","111100","111101","111100","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","101000","101001","100101","010101","010101","010110","010101","010101","010101","101001","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","101001","101001","010101","010101","010110","000110","010110","000110","000101","101001","111001","111101","111100","111100","111100","111100","111100","111100","111100","111100","101000","101001","010101","010101","010101","101001","111101","111100","111100","111100","111100","111100","111000","101000","010100","111000","111100","111100","111000","101001","010101","010110","010110","010101","101001","111101","111100","111100","111100","111100","111000","111000","101000","101001","010101","010101","010110","010110","000110","000110","000110","000110","000110","000110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111000","101000","101001","010101","010110","010101","010100","111001","111100","111100","111000","111000","111000","111100","111100","111100","111100","111100","111000","101000","101000","101000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010110","000110","010110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000001","000101","000101","000001","000110","000110","010110","010110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","111101","111100","111100","111100","111100","111100","111101","111001","101001","010101","010110","010110","000110","000110","000110","010110","010101","111001","111100","111100","111100","111100","111100","111000","101000","101001","010101","010101","000110","010110","000110","000110","000110","010101","010101","010101","010101","010101","010101","010110","010101","010100","111001","111100","111100","111100","111000","111000","101001","010101","000110","010110","010101","101001","111100","111100","111100","111100","111100","111100","101000","101000","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","101001","101001","010101","010101","010101","010110","010110","010101","010101","101001","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","101001","101001","010101","010101","010110","010110","010110","000110","010110","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","010101","010101","010101","010101","010100","111101","111100","111100","111100","111100","111100","101000","010100","010100","111001","111100","111100","111000","101001","010101","010101","010110","010101","101001","111101","111100","111100","111100","111100","111100","111000","111000","101000","101001","100101","010101","010110","000110","000110","000110","000110","010110","010110","010110","010101","100101","101001","111101","111100","111100","111100","111100","111000","101000","100101","010101","010110","010101","010100","111001","111100","111100","111000","101000","101000","111100","111100","111100","111100","111100","111000","111000","111000","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","100101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000101","000101","000110","000110","000110","010110","000110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111100","111100","111100","111100","111100","111100","111100","111001","101001","010101","010101","010110","010110","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111000","111000","111001","100101","010101","010110","010110","000110","010110","000110","000110","000110","000110","000101","010110","010110","010110","010101","101000","111101","111100","111100","111100","111000","101000","101001","010101","000110","010110","010101","101001","111100","111100","111100","111100","111100","111000","010100","010100","101001","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111100","111000","111000","101000","101001","010101","000101","000110","010110","010110","010101","010101","010101","101001","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111001","111001","101001","101001","010101","010101","010101","010110","000110","000110","000110","000110","010110","010101","010101","101000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","010101","010110","000110","010110","010100","101001","111100","111100","111100","111100","111000","101000","010101","010100","101001","111101","111100","101000","101001","010101","010101","010101","010101","101001","111101","111100","111100","111100","111100","111100","111000","111000","101000","101000","101001","100101","010101","010101","010101","010110","010110","010110","010101","010101","100101","111001","111100","111100","111100","111100","111100","111100","111000","101001","010101","010101","010110","000101","010100","111101","111100","111000","111000","100100","101000","111100","111100","111100","111100","111100","111100","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010101","000110","010110","000110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000001","000101","000110","000001","000110","000110","000110","010110","010110","010101","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","010101","010101","010110","000110","000110","000110","000110","000110","010101","101001","111101","111100","111100","111100","111100","111100","111000","111000","101000","101001","010101","010101","010110","000110","000110","000110","000110","000110","010110","010110","000110","000110","010101","010101","101000","111100","111100","111100","111100","111100","101000","101001","010101","000110","010110","010101","111001","111100","111100","111100","111100","101000","101000","010100","010101","010101","010100","101001","101001","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","101000","101001","010101","010101","000110","000110","010110","010110","010101","010101","010101","101001","111001","111101","111100","111100","111100","111101","111101","111101","111101","111101","111101","111101","111001","101001","101001","010101","010101","010101","010110","010110","010110","000110","000110","000110","010110","010110","000110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010110","010110","010110","010101","010100","111101","111100","111100","111100","101001","100101","010101","010101","100101","111101","111000","101000","101001","010101","010101","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111000","111000","101000","101000","101001","101001","100101","010101","010101","010101","010101","100101","101001","111001","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010101","000110","010101","101000","111101","111100","111000","111000","100100","101000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000001","000101","000101","000101","000101","000110","010110","010110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111001","101001","010101","010101","000101","010110","010110","000110","000110","000110","000110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","101001","010101","010101","010110","000110","000110","000110","010110","000110","000110","000110","010110","010101","101001","111100","111100","111100","111100","111100","111000","101000","101001","010101","000110","010110","010101","111001","111100","111100","111100","111100","101000","101001","010101","010101","010101","010101","010101","010101","100101","111001","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","101000","101001","010101","010101","010110","010110","010110","010110","010101","010101","010101","010101","010101","101001","101001","101001","101001","101001","101001","101001","101001","100101","010101","010101","010101","010101","010101","010110","010110","010110","010110","000110","010110","010110","010110","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","101001","010101","010110","000110","000110","010101","010100","101001","111101","111100","111000","101001","010101","010101","010101","010100","111101","111000","101000","101001","010101","010101","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","111000","111000","101000","101000","101000","101000","101000","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","101001","010101","010110","000101","010101","101001","111100","111100","111000","101000","010100","101000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","100101","010101","010110","000110","000110","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000101","000001","000101","000101","000101","000110","000110","000110","000110","000101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111001","101001","010101","010101","010110","000110","000110","000110","000110","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","101001","101001","010101","010101","010101","010101","000101","000101","010101","010110","010101","010101","101001","111001","111100","111100","111100","111100","111100","111000","101001","100101","010101","010110","010110","010101","111001","111100","111100","111100","111100","101000","101001","010100","010101","010110","010110","010110","010110","010101","010101","101001","111001","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","101000","101001","010101","010101","010101","000110","010110","010110","010110","010110","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010110","010110","010110","010110","010110","010110","010110","000110","000110","010110","010110","000110","000110","010110","010110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","101001","010101","010110","000110","000110","010110","010101","010100","111101","111101","111001","101001","010101","000110","010101","010101","111101","111001","101000","101001","010101","010101","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","111000","111000","111000","111000","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010101","000101","010110","010101","010100","111101","111100","111101","111000","101001","010100","101000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010110","000110","000110","000110","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","000001","000101","000001","000101","000001","000110","000110","000110","000110","000110","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111001","100100","010101","010101","000110","000110","000110","000110","000110","000110","000110","000110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","101000","101001","101001","010101","010101","010101","010101","010101","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111000","101001","010101","010101","010110","010101","010101","111101","111100","111100","111100","111100","101000","101001","010101","010101","010110","010110","010110","010110","010110","010110","010101","010101","010101","111001","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","111000","101001","010101","010101","010101","010101","010110","010110","010110","010110","010110","000110","010110","010110","000101","010110","010110","010110","010110","010110","000110","000110","000110","000110","000110","000110","010110","010110","010110","000110","000110","000010","000010","010110","010110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010110","000110","000110","010110","000101","010101","101001","111101","101001","010101","010101","010110","000101","010101","111001","111001","101000","101001","010101","010101","010101","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111001","101001","010101","000101","010110","010101","101001","111101","111100","111100","111000","101001","010100","101000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000001","000001","000001","000001","000110","000110","000110","000110","000110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010101","010110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","101000","101000","101001","101001","101001","101001","101001","101001","111001","111101","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010110","010110","010101","010101","111101","111100","111100","111100","111100","101000","101001","010101","010101","010110","010110","010110","010110","010110","010110","010110","010110","010101","010101","101001","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","101000","111001","101001","010101","010101","010101","010101","010101","010110","010110","000110","010110","010110","010110","000110","010110","010110","010110","010110","000110","000110","000110","010110","010110","010110","000001","000110","000101","000001","000001","000001","000110","010110","010110","010101","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111001","100101","010101","000110","000110","000110","000110","000110","010101","010101","101010","101001","010101","000110","010110","000101","010101","101001","111001","101000","101001","010101","010101","010101","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111100","111101","101001","010101","010101","010110","010101","010101","101001","111100","111100","111000","101000","101001","010100","101000","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","100101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000001","000101","000001","000001","000010","000110","000110","000110","000110","010110","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010101","000110","000110","000110","000110","000110","000101","000101","000110","010110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","111000","111000","101000","101000","101000","111000","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","100101","010101","010110","010101","010101","101001","111100","111100","111100","111100","111100","101000","101001","010101","010101","010110","010110","010110","000110","000110","000110","000110","000110","010110","010110","010101","010101","101001","101001","111101","111101","111100","111000","111100","111100","111100","111100","111000","111000","111000","111000","111000","101000","101001","101001","100101","010101","010101","010101","010101","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","000110","000001","000001","010110","011010","000101","000001","000001","000001","010110","010110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010101","000110","000110","000110","000110","000110","010110","010101","101010","010101","010110","010110","010110","000101","010101","101001","111001","101000","101001","100101","010101","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111101","111001","010101","010101","010110","010101","010101","101001","111101","111100","111100","111000","101000","010101","010100","101000","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010101","010110","010110","000110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000101","000001","000001","000001","000110","010110","000110","000110","010110","010101","101001","111101","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010110","000110","000110","000110","000110","000110","000101","000101","000110","010110","010110","010101","010101","111001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","111000","111000","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","010101","010101","010110","010101","010101","111101","111100","111100","111100","111100","111100","101000","101001","010101","010101","010110","010110","010110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010101","010101","100101","101001","111101","111101","111100","111100","111100","111100","111100","111100","111000","111000","111000","111000","111000","101000","101000","101001","101001","100101","010110","010110","010110","010110","000110","000110","000110","000110","000110","000110","000110","000001","000001","010110","010110","101111","101111","000001","000001","000001","000001","010110","010110","010110","010110","010101","101001","111101","111101","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010101","000110","010110","010110","000110","010110","010110","000110","010110","010110","010110","010110","010110","000110","010101","101001","111101","111000","111000","101001","010101","010110","010110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111001","101001","010101","000101","010101","010101","010100","111001","111101","111100","111100","111000","101001","010101","010100","101000","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000001","000001","000001","000001","000001","010110","000110","010110","010110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101001","010101","010101","000110","000110","000110","000110","000110","000101","000101","000110","000110","000110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010110","000101","010101","010100","111101","111100","111100","111100","111100","111100","101000","101001","010101","010110","010110","000110","000110","000101","000101","000110","000110","000110","000110","000110","000110","010110","010110","010101","010101","010101","100101","111001","111101","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","111000","111000","101000","101000","101001","101001","010110","010110","010110","010110","000110","000101","000001","000001","000001","000001","010101","101010","000000","000000","000000","101011","000001","000001","000001","000001","010110","010110","010110","010110","010110","101010","101010","111001","111001","111101","111101","111101","111100","111101","111101","101001","101001","010101","010101","000110","010110","010110","000110","000110","000110","000110","010110","010110","010110","010110","010110","010110","010101","011001","111101","111000","111000","101001","010101","010101","000110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","010101","010101","010101","010101","101001","111101","111100","111100","111100","111000","101001","010101","010101","101000","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","101001","010101","010110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000001","000001","000101","000001","000101","010110","010110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","101001","010101","000110","000110","000110","000110","000110","000101","000101","000110","000110","000110","000110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010101","010101","000110","010101","010101","101001","111101","111100","111100","111100","111100","111100","101000","101001","010101","010101","010110","000110","000110","000001","000001","000101","000110","000101","000110","010110","000110","000110","000110","010110","010110","010110","010101","010101","101001","111001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","111000","101000","101001","010101","010101","010110","000110","000110","000110","000101","010101","101010","000000","000000","000000","000000","000000","000000","101010","000001","000001","000001","000001","010110","010110","010110","000110","000101","010110","010101","010101","010101","010101","101001","101001","101001","111101","111101","101001","101001","010101","000101","010110","010110","010110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010110","010101","111101","111000","111000","101000","101001","010101","000101","010110","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","101001","010101","010101","010110","010101","010101","101001","111101","111100","111100","111100","111100","111000","101001","010101","010101","101000","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","010101","010101","010110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000001","000001","000101","000001","000001","000110","000110","010110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010110","000110","000110","000110","000110","000101","000101","000110","000110","000110","000110","010101","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111001","100101","010101","010110","010110","010101","010101","111101","111100","111100","111100","111000","111100","111100","111000","101001","010101","010101","000110","000110","000110","000110","000001","000110","000001","000101","000101","000110","000110","000110","000110","000110","000110","010110","010110","000101","010101","010101","101001","111001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","100101","010101","010110","010110","010110","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","010101","000001","000001","000001","000110","000110","010110","000110","000110","000110","000110","010110","010101","010101","010101","010101","010101","010101","010101","010101","010101","010110","010110","000110","010110","010110","000010","000110","000110","000110","000110","000110","000110","010110","000110","010110","010110","010110","010101","111101","111100","111000","101000","101000","010101","010101","010110","010110","010101","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111001","101001","010101","010101","000101","010101","010101","100101","111001","111101","111100","111100","111100","111100","101000","101001","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010101","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","000001","000001","000001","000101","000001","000101","010110","010110","010110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010110","000110","010110","000110","000110","000101","000101","000110","000110","000110","000110","010110","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","010110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","101000","101001","010101","010101","000110","000110","000110","000110","000001","000101","000001","000001","000101","000001","000101","000110","000110","000110","000110","000110","000110","010110","010110","010101","010101","010101","101001","111001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","100101","010101","010110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000001","000001","000001","000001","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010110","010101","010101","010110","010110","000110","000110","000110","000010","000010","010110","000110","000110","000110","010110","000110","010110","000110","010110","010110","010110","010101","111101","111101","111000","101000","111000","101001","010101","010110","010110","010110","010101","010101","111001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","101001","010101","010101","010110","010110","010101","010100","111001","111101","111100","111100","111100","111100","111100","101000","101001","010101","010101","100101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010101","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000001","000001","000101","000001","000001","000110","010110","000110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010101","010110","010110","000110","000110","000101","000101","000110","000110","000110","000110","010110","010101","101001","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","010101","010110","010110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","101000","101001","010101","010101","000110","000110","011010","000000","011010","000001","000001","000101","000001","000001","000001","000001","000110","000110","000110","000110","010110","010110","010110","010110","010110","010101","010101","010101","101001","111101","111101","111100","111100","111100","111100","111100","111100","111000","101000","100101","010101","010110","000110","000110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000001","000001","000001","000001","000110","000110","000110","010110","000110","000110","000110","000110","000110","010110","000110","000110","010110","010110","010110","000110","010110","000110","000110","000110","000110","000010","000010","000010","000110","010110","000110","010110","010110","000110","000110","010110","010110","010110","010101","101001","111100","111000","111000","111000","101001","101001","010101","010101","010110","010110","010101","010101","101001","111101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","101001","011001","010101","010101","010110","010110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111000","101000","100101","010101","010101","100101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010101","010110","010110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000001","000101","000001","000001","000001","000101","010110","000110","010110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","100101","010101","010110","010110","000110","000110","000110","000001","000101","000110","000110","000110","010110","010101","010101","101001","111101","111100","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","010101","000110","010110","010110","010110","010101","111001","111100","111100","111100","111100","111100","111100","111100","101000","101001","010101","010101","000110","010110","010110","000000","000000","000000","011010","000101","000001","000001","000001","000001","000001","000001","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010101","010101","101001","111001","111101","111100","111100","111100","111100","111000","101000","100101","010101","010110","010110","000110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000001","000001","000001","000101","000001","000001","000001","000001","000001","000101","000110","010110","010110","010110","010110","010110","000110","000110","000110","010110","000110","000110","000110","010110","000110","000110","000001","000010","000110","000110","000110","010110","010110","000110","000110","010110","010110","000110","010101","101001","111101","111100","111000","111000","111000","101001","101001","010101","010101","010110","010110","000101","010101","010101","101001","111001","111101","111101","111101","111101","111101","111101","111101","111001","101001","101001","010101","010101","010110","000110","000110","000110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111000","101001","010101","010101","010101","100101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010101","000001","000001","000001","000001","000001","000110","000110","010110","010110","010101","100100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010110","010110","000110","000110","000110","000001","000110","000110","000110","010110","000110","010110","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","010101","010110","010110","000110","010110","010110","010101","111001","111100","111100","111100","111100","111100","111100","111100","101000","101001","010101","010101","010110","000110","011010","000000","000000","000000","000000","000000","101010","000001","000001","000101","000101","000001","000001","000001","000101","000110","010110","010110","000110","000110","000110","000110","010110","010101","010101","010101","100101","111001","111101","111101","111100","111000","101000","100101","010101","010110","010110","000110","101011","000000","000000","000000","000000","000000","000000","000000","000000","101011","010101","000001","000001","000001","000001","000101","000101","000001","000001","000001","000001","000001","000001","000001","000101","000110","000110","000101","000110","000110","010110","000110","010110","000110","010110","000001","000001","000101","000101","000110","000110","010110","000110","000110","000110","010110","010110","000110","010101","101001","111101","111100","111100","111000","111000","111000","101001","100101","010101","010101","010110","010101","010101","010101","010101","010101","010101","010101","100101","100101","100101","010101","010101","010101","010101","010101","010101","010110","010110","010110","010110","000110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010101","010101","100101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","010101","010101","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","000001","000001","000001","000001","000001","000101","010110","010110","010110","010101","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010110","010110","000110","000110","000110","000010","000110","000101","000001","000110","000110","010110","010110","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","101001","010101","010101","010110","010110","000110","000110","010110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","011010","000001","000001","000101","000001","000001","000101","000001","000001","000110","000110","000110","000110","010110","010110","010110","010110","010101","010101","010101","101001","101001","111101","101001","101001","010101","010101","010110","000110","000110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","101011","011010","010110","000001","000001","000001","000001","000001","000101","000001","000001","000001","000001","000001","000001","000101","000101","000001","000001","000101","000110","000110","000001","000001","000101","000001","000110","000110","010110","000110","000001","000110","010110","010110","000110","010101","010100","111101","111100","111000","111000","111000","111000","111000","101001","101001","010101","010101","010101","010110","010110","010110","010101","010101","010101","010101","010101","010110","010101","010110","010101","010110","010110","010110","010110","000110","000110","000110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","101000","101001","010101","010101","010101","100101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","010101","010110","010110","010110","000110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000001","000001","000001","000001","000001","000001","010110","010110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101000","010101","010101","010110","000110","000110","000110","000010","000001","000110","000001","000101","010110","000110","010110","010110","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111001","101001","010101","010101","000110","010110","000110","000110","000110","010110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","101000","101001","010101","010101","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000001","000001","000001","000001","000001","000001","000001","000101","000110","000110","010110","000110","000110","010110","010110","010110","010101","010101","010101","101001","101001","101001","011010","010110","010110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","101011","011010","010101","000101","000001","000001","000001","000001","000001","000001","000001","000001","010101","010110","101011","000101","000101","000001","000001","000101","000001","010110","000110","000101","000001","000110","000110","010110","010110","010101","010100","111101","111101","111100","111100","111000","111000","111000","101000","101000","101000","011001","010101","010101","010110","000110","010110","010110","010110","000110","000110","000110","000110","000110","010110","000110","000110","010110","000110","000110","010110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","101000","101001","010101","000110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010110","010110","010110","000101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000001","000001","000001","000001","000001","000110","010110","000110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","000110","010110","000110","000110","000110","000001","000001","000001","000101","000110","010110","000110","000110","010110","010101","010101","101001","111001","111101","111101","111100","111100","111100","111100","111100","111000","111100","111101","111101","111101","111001","101001","010101","010101","010110","010110","000110","000110","000110","000110","000110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111101","101001","101001","010101","010110","010110","000110","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000101","000001","000001","000001","000001","000001","000001","000001","000110","000110","000110","000110","000110","000110","010110","010110","010101","010101","010101","010101","010110","010110","010110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","101010","010101","000001","000001","010101","101010","000000","000000","010110","000101","000001","000001","000101","000001","000110","000101","000001","000001","000010","000110","000110","000110","010101","010101","101001","111101","111101","111101","111101","111100","111000","111000","101000","101000","101001","101001","010101","010101","010110","010110","010110","010110","010110","000110","000110","010110","000110","000110","010110","000110","000110","000110","000001","000110","000110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","101000","010101","010110","000110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","100101","010101","010110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000001","000001","000001","000001","000001","000110","000110","000110","000110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","000110","010110","000110","010110","010110","000110","000001","000101","000001","000001","000110","000110","000110","010110","010110","010101","010101","010101","100101","101001","111001","111101","111101","111101","111101","111101","111101","101001","101001","010101","010101","010101","010101","010110","010110","000110","000110","000110","000110","000110","000110","000110","010110","010101","101001","111101","111101","111100","111101","111101","111101","111101","101001","101010","010101","010110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000001","000001","000001","000001","000001","000001","000001","000101","000101","000110","000110","010110","000110","000110","010110","010110","010101","010101","010110","000110","010110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000001","000001","000001","000101","000001","000001","000001","000001","000001","000110","000110","000110","000110","000101","010101","101001","101001","101001","101001","111001","111101","111001","111001","101001","101001","101010","010110","010110","000110","000110","000110","000110","000110","000110","000110","000110","010110","000101","000101","000001","000001","000001","000001","010110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111000","101000","010101","010110","010110","010101","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","010101","010101","010110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010101","000001","000001","000001","000001","000001","000110","010110","000110","000110","010101","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010101","010110","000110","010110","011011","010110","000001","000010","000001","000010","000001","000110","010110","000110","000110","010110","010110","010110","010101","010101","010101","010101","010100","010101","011001","010100","010100","010101","010101","010101","010110","010110","010110","010110","000110","000110","000110","000110","000101","000101","000110","010110","010110","010101","010110","111010","101001","101001","101001","101001","010101","010101","010101","010101","000101","000110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000001","000001","000001","000001","000001","000001","000101","000101","000101","000110","000110","010110","010110","000110","010110","010110","010110","000110","000110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000001","000001","000001","000001","000001","000001","000001","000001","000001","000110","000110","000110","000110","010110","010101","000101","010101","010101","010101","010101","010101","100101","101001","101001","101001","101010","010110","010110","010110","010110","000110","000110","000101","000001","000001","000101","010110","101011","011010","000001","000001","000001","000010","010110","010110","010110","010101","101010","111101","111101","111100","111100","111100","111100","111100","111000","101001","010101","010110","010110","010101","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010101","010110","010110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000001","000001","000001","000001","000001","000101","010110","000110","010110","000110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101001","101001","010101","010110","000110","010110","010110","000000","010110","000001","000010","000001","000001","000001","000101","000110","000110","000110","010110","000110","000110","010110","010110","010101","010101","010101","010101","010101","010101","010110","010110","000110","000110","000110","000110","000110","010110","000110","000110","000110","000101","000110","000110","000110","010110","010110","010110","010101","010101","010101","010101","010101","010101","010101","010101","010110","000110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000001","000001","000101","000001","000001","000001","000001","000101","000110","000110","000110","010110","000110","000110","010110","010110","000110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000001","000001","000101","000001","000001","000001","000001","000001","000001","000110","010110","010110","000110","010110","000110","000110","000110","000110","010110","010101","010101","010101","010101","010101","010101","010110","010110","010110","010110","010110","000110","000110","011010","101010","101111","000000","000000","000000","010110","000001","000001","000001","000010","010110","000110","000110","010110","101010","101001","111101","111101","111101","111101","111101","111101","111001","101001","010101","010110","000110","010101","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","100101","010101","010110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010101","000001","000001","000001","000001","000001","010110","000110","000110","000110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010110","010110","010110","010110","000000","101011","010110","000001","000001","000101","000101","000001","000101","000110","010110","000110","000110","010110","010110","000110","000110","000110","000110","000110","010110","010110","000110","000110","010110","000110","000110","000110","000101","011010","010110","000101","000101","000110","000110","000110","010110","010110","010110","000110","000110","000101","010101","010110","000101","010110","010110","000110","000110","000110","010110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000101","000001","000001","000001","000001","000001","000010","000110","000110","000110","000110","000110","000110","000110","000110","010110","000110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","000101","010110","000000","010110","000001","000001","000001","000001","000110","010110","010110","010110","010110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010110","010110","010110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","010101","000001","000001","000001","000110","000110","000110","010110","010110","010101","010101","010100","010100","100101","101001","101001","101001","101001","100101","010110","010110","000110","010101","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010101","010101","010110","010110","010101","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","000001","000001","000001","000001","000001","000110","010110","000110","000110","010110","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","000110","010110","010110","000110","101011","000000","101011","010101","000001","000001","000001","000001","000001","000001","000001","000110","000110","000110","000110","000110","010110","010110","010110","010110","000110","010110","010110","010110","000110","000110","000110","000101","101011","000000","011010","000101","000110","000110","000110","000110","000110","000110","000110","010111","000110","000110","000110","000110","010110","010110","010110","000110","000110","010110","000110","000110","010101","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000001","000001","000001","000001","000001","000001","000001","000001","000101","000101","000110","000110","010110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000001","000001","000001","000001","000001","000110","010110","000110","010110","010110","010110","000110","000110","000110","000110","000110","000110","000110","010110","000110","000110","010110","000110","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","010001","000001","000001","000001","000110","000110","000110","000110","000110","000110","010101","010101","010101","010101","010101","010101","010101","010101","010101","010110","010110","000110","000101","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010110","000110","010110","010101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000001","000001","000001","000001","000001","010110","000110","000110","010110","010101","100101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010101","000110","010110","010110","011010","000000","000000","000000","000101","000101","000001","000001","000001","000001","000001","000001","000101","000101","000110","000110","000110","010110","010110","010110","010110","010110","010110","000101","000001","000001","010101","101111","000000","000000","011010","000101","000110","000110","000001","000110","010110","010110","010110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","000110","000101","000101","101010","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000001","000001","000001","000001","000001","000001","000001","000101","000101","000110","010110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000110","000110","010110","000110","000110","000110","000110","000110","000110","010110","000110","000110","000110","000110","000110","010110","000101","000000","000000","000000","000000","000000","000000","000001","000001","000001","000001","000110","000110","000110","000110","000110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","000110","010101","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111001","100101","010101","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","000001","000001","000001","000001","000001","000110","010110","000110","010110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111000","111000","101001","010101","010101","010110","010110","010110","010110","000000","000000","000000","000000","011010","000001","000001","000001","000001","000001","000101","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000101","101010","000000","000000","000000","000000","011010","000110","000110","000001","000110","010110","000110","000110","010110","000110","010110","000110","000110","000110","000101","000110","000110","000001","000001","000001","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000001","000001","000001","000001","000001","000001","000001","000001","000110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010101","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000101","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","101111","000000","000000","000000","000000","000000","000001","000001","000001","000001","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","000110","000110","000110","000110","010101","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010101","000110","010110","000101","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000001","000001","000001","000001","000001","000001","010110","000110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","010110","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","010101","101010","000000","000000","000000","000000","000000","000000","101011","010110","000110","000110","000001","000001","000110","000101","000001","000001","000001","000001","000001","000001","000001","000001","000001","010110","101010","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000001","000001","000001","000001","000001","000001","000001","000001","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","011010","010101","000101","000000","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000110","000110","010110","000110","010110","101011","000000","000000","000000","000000","111011","000001","000001","000001","000001","000001","000001","000001","000001","000101","000101","000110","000110","000110","000110","000110","000110","000110","010110","000110","000110","000110","000110","000101","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000001","000001","000001","000001","000001","000110","010110","000110","010110","010101","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","000110","010110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","101011","010101","000101","000001","000001","000001","000001","000001","000001","000101","000101","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","000001","000001","000101","000001","000001","000001","000001","000001","000001","010110","010110","101010","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000001","000001","000000","000001","000101","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","101010","010101","010101","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","010110","101011","000000","000000","000000","000000","101010","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000101","000101","000110","000110","000110","010110","010110","010110","010101","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111000","100101","010101","010110","000110","000110","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000001","000001","000001","000001","000001","000001","010110","000110","010110","010110","010101","101001","111101","111000","111100","111100","111100","111100","111100","111100","111000","101000","101001","010101","010110","010110","010110","000110","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","010101","010101","010110","101010","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000101","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","100110","010110","000001","000001","000001","000001","000001","000001","000001","000001","101011","000000","000000","000000","000000","000000","000000","000000","101011","101011","101010","010110","010101","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000110","000110","010110","010101","010101","111101","111101","111100","111100","111100","111100","111100","111100","111100","101001","010101","010110","010110","010110","000101","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010101","000001","000001","000001","000001","000001","000110","000110","000110","010110","010101","010101","111001","111100","111100","111100","111100","111100","111100","111100","111000","111001","101001","011010","000110","010110","010110","010110","010101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","010110","010101","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","101010","010110","010101","000001","000001","000001","000001","000001","000001","000001","000110","000110","010110","010110","010101","111101","111101","111100","111100","111100","111100","111100","111100","111000","101001","010101","010110","010110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","000001","000001","000001","000001","000001","000110","000110","000110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111101","111001","101001","100101","010101","000110","000110","000110","010110","010101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000001","000001","000001","000001","000110","010110","010110","010110","010101","101001","111101","111101","111101","111100","111100","111100","111100","101000","100101","010101","010110","010110","000110","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000001","000001","000001","000001","000001","000110","000110","010110","010110","010101","101001","111101","111101","111101","111101","111101","101001","101001","010101","010101","010101","010110","000110","010110","010110","010110","010101","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000001","000001","000001","000001","000101","000110","010110","000110","010110","010101","010101","100101","101001","111001","111101","111101","111101","101001","010101","010101","010110","010110","000110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","000001","000001","000001","000001","000001","000101","010110","000110","010110","010101","010101","101010","101001","101001","101001","010101","010101","010101","010101","010110","000101","010110","000110","000110","010110","010110","010101","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000001","000001","000001","000001","000001","010110","010110","000110","010110","010110","010101","010101","010101","010101","100101","101001","101001","101001","010101","010110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000001","000001","000001","000001","000001","000001","000110","010110","010110","000110","010110","010110","010101","010101","010101","010110","010110","010110","000110","010110","010110","000110","010111","010110","000110","010110","010101","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000001","000001","000001","000001","000001","010110","010110","010110","010110","010110","010110","010110","010101","010101","010101","010101","010101","010101","010110","010110","010110","010110","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000000","000001","000001","000001","000001","000101","000110","010110","000110","000110","010110","000110","010110","010110","000110","000110","010110","010110","010110","000110","010110","000110","010110","010110","010101","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000001","000001","000001","000001","000001","000101","000110","010110","000110","000110","000110","010110","010110","010110","010110","000110","000110","000110","000110","010110","010110","010110","101011","000000","000000","000000","000000","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000001","000001","000001","000001","000001","000001","000110","000110","000110","010110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000001","010101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000001","000001","000001","000001","000001","000001","000001","000001","000110","000110","000110","000110","000110","000110","000110","000110","010110","000110","000110","000110","000110","010110","000000","000000","000000","000000","101010","101010","010101","000000","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000000","000001","000001","000001","000001","000110","010110","000110","000110","000110","010110","000110","000110","000110","000110","010110","000110","000101","000001","000001","000001","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010101","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000101","000110","010110","000110","000110","000110","000110","000110","000110","010110","010110","000000","000000","000000","000000","101010","101010","101011","000000","010101","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000001","000001","000001","000001","000001","000010","000110","010110","000110","000110","000110","010110","000110","000101","000001","000001","000001","010101","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","010110","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000101","000110","000110","010110","000110","010110","010110","101011","000000","010101","000000","000000","010101","101010","101010","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000000","000001","000001","000001","000001","000110","010110","010110","000110","000110","000001","000001","000001","010101","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","010110","000001","000001","000001","000001","000001","000001","000001","000001","000001","000001","000101","000101","000101","010110","000000","000000","000000","000000","111110","010101","000000","101011","010101","000000","010101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","000000","000101","000001","000001","000001","000001","000101","000001","000001","000001","010101","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","010110","010001","000001","000001","000001","000001","000001","000001","000001","000001","010101","101011","000000","000000","010101","000000","000000","000000","010101","010101","000000","000000","010101","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000001","000000","000001","000001","000001","000001","000001","010101","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111011","100110","010001","000001","000001","000001","000101","101010","000000","000000","000000","000000","000000","000000","000000","010101","000000","010101","000000","000000","010101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000001","000001","000001","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","101010","101010","000000","000000","000000","000000","000000","000000","101010","101010","000000","010101","000000","101010","010101","000000","010101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010101","101010","000000","000000","000000","101010","010101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","011010","010110","010110","010110","010110","010110","010110","010110","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","011010","010110","010110","010110","010110","010110","010110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","010110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","011010","010110","010110","010110","000110","010110","010110","000110","010110","010110","000110","010111","000110","000110","000110","000110","010110","000110","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","011010","010110","010110","010110","000110","000110","000110","000110","010110","010110","010110","000110","000110","000110","000110","010110","010110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","010110","010110","010110","000110","000110","010110","010110","010110","010110","000110","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","101011","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","011010","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","010110","010110","010110","010110","010110","010110","000110","000110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","000110","000110","000110","000110","000110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","101011","010110","010110","010110","010110","010110","000110","010110","000110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","000110","010110","000110","000110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","010110","010110","010110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","010110","010110","010110","000110","010110","010110","000110","010110","010110","010110","000110","000110","000110","000110","000110","000110","010110","010110","000110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","101011","010110","010110","010110","010110","000110","000110","000110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010101","010101","010110","010110","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","011010","010110","010110","010110","010110","010110","010110","010110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010110","010101","010101","000110","000110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","010110","010110","010110","000110","000110","000110","010111","000110","000110","010110","010110","010110","010110","010110","010110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","010110","010110","010110","000110","000110","010110","000110","000110","000110","000110","010110","000110","010110","010110","010110","010110","010110","000110","000110","000110","010110","000110","000110","000110","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","010110","010110","000110","000110","010110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010110","010110","010110","010110","010101","010101","010101","010101","010101","010101","010101","101001","101010","101110","111110","101010","010110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","010110","000110","010110","000110","000110","000110","010110","000110","000110","000110","000110","000110","000110","010110","010110","000110","000110","010110","010110","010110","010110","010110","010101","010101","010101","010101","010101","010101","010101","101001","111010","111110","101010","011010","010110","000110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","010110","010110","010110","010110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010101","010101","011001","101010","101010","010110","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","011010","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","010110","010110","010110","000110","010110","010110","000110","000110","000110","000110","010110","000110","010110","010110","010110","010110","010110","010101","010101","010101","010101","010101","010101","010110","010110","010110","010110","000110","000110","000110","000110","010110","010110","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","010110","010110","000110","000110","000110","000110","000110","000110","010110","010110","000110","000110","000110","010110","010110","010110","010110","010101","010101","010101","010101","010100","010100","101001","101001","111101","111101","111101","111101","111101","111101","111100","111100","111100","111101","101001","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","010110","010110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","000110","010110","010110","010101","010101","010101","010101","010100","010100","101001","101001","111001","111101","111101","111101","111101","111101","111101","111100","111100","111100","111101","101001","010101","000110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","010110","000110","000110","000110","000110","000110","000110","010110","010110","010101","010101","010101","010100","111001","111101","111101","111101","111101","111110","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010101","010101","010101","010101","010101","101001","101001","101001","111101","111101","111101","111001","101001","101001","010101","010101","010101","010110","010110","000110","000110","000110","000110","000110","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","000110","000110","000110","000110","010110","010110","010110","010110","010110","010101","010101","010101","010101","010101","010101","011001","101001","111110","111101","111101","111101","111101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010101","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","000110","010110","010110","010110","010110","010110","010110","010101","010101","010101","010101","010101","010101","010101","101001","101110","111110","111101","111101","111101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","000110","000110","000110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","010110","000110","000110","010110","000110","010110","010110","010101","010101","010101","101001","111110","111101","111101","111100","111100","111100","111100","111100","111101","010101","010110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","010110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000110","010110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010101","010101","010101","011001","101001","111110","111101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111101","111101","111101","111101","111101","101001","010101","010110","010110","010110","000110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","000110","010110","010101","010101","010100","010100","101001","111001","111101","111101","111101","111101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010110","010101","010101","010100","010100","101001","111101","111101","111101","111101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111110","010101","010110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","010110","000110","000110","010110","010110","010101","010101","101001","111101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","010110","010110","010110","010110","000110","000110","000110","000110","010110","010110","010110","010101","010101","010101","010101","010101","010110","010110","010110","000110","000110","000110","000110","000110","010110","010110","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","010110","000110","000110","000110","000110","010110","010110","010110","010101","010101","010100","101001","111101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","010110","000110","010111","010110","000110","010110","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010101","111110","111101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","000110","000110","010110","101010","111110","111101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111110","010101","010110","000110","010110","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","000110","010110","010110","101001","111110","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","000110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000110","010110","000110","010111","000110","010110","010110","010101","010101","010101","010101","101001","101001","101010","111110","111110","101001","101001","011001","010101","010101","010101","010110","010110","010110","000110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","000110","010110","010110","010101","010101","010101","101001","111101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","010101","010110","000110","000110","010110","010110","101111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","010110","000110","010110","010110","101010","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111110","010101","010110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111110","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000110","000110","000110","000110","000110","010110","010101","010101","101001","111101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","101001","010101","010110","000110","010110","000110","000110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","010110","000110","010110","010101","011001","101001","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000110","000110","000110","010101","111110","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","010110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","010110","010101","010101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","101001","010101","010110","000110","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","000111","010110","011001","111110","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","010110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","010110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000110","000110","000110","010101","111110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","010111","010110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","000110","010110","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000110","000110","000110","000110","010110","010101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","011001","010110","010110","000110","000110","010110","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000110","000110","000110","010110","010101","111110","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111001","010101","010110","000110","000110","000110","101111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010110","000110","000110","000110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000110","000110","000110","000110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010101","101010","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010110","000110","000110","000110","101011","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","010110","010110","010101","111110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111110","010101","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000111","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000110","000110","000110","010110","010110","101001","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010110","000110","000110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010110","000110","000110","010110","101011","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","111101","111101","111110","011010","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","010110","010110","010101","111110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","111101","111101","111101","101110","010101","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","111110","111101","111101","111101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010110","100100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010110","000110","000110","010110","101011","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","111101","111101","111101","111101","111110","111110","101101","101001","101001","010101","010101","010101","010101","010110","010110","000110","000110","000110","000110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","111101","111101","111101","111101","111101","111110","111110","101001","101001","010101","010101","010101","010101","010101","010110","000110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000111","000110","010110","010101","010101","010101","010101","010101","101000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","000110","000110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","010110","000110","010110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","010110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","111101","111101","111101","111101","111110","111110","111001","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","011001","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","010100","010100","010100","010101","010101","010101","010101","010101","010101","010101","010110","010110","010110","000110","010110","000110","000110","000110","000110","000110","101011","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","100100","010100","010100","010101","010101","010101","010101","010101","010101","010101","010110","010110","010110","000110","000110","000110","000110","000110","000110","000110","010110","000000","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","101000","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","010110","011001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","000110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111101","111101","101001","010100","010100","010101","010101","010101","010101","010101","010101","010100","101000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010101","000110","000110","000110","000110","101111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","010110","010110","101010","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","010110","010110","010110","010110","010110","010110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","000110","000110","000110","010110","010101","111110","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","010101","010110","010110","010110","010110","010110","010110","010110","010110","000110","000110","000110","000110","000110","010111","000110","000110","000110","000110","000110","000110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","000110","000110","000110","000110","010110","000110","000110","000110","010110","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010101","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111101","111101","111010","010101","010101","010101","010110","010110","010110","010110","010110","010110","010110","010101","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","010110","000110","010110","010110","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","101010","111110","111101","101000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","000111","000110","000110","000110","010110","000110","000110","000110","000110","010110","010110","010110","010110","010110","010110","000110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","000110","000110","010110","010101","101110","111110","111101","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010110","010110","010110","010110","000110","000110","010110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","010110","010110","000110","000110","010110","010110","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","010110","000110","000110","010110","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","000110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","101001","111101","111100","111101","111101","101001","010101","010101","010110","010110","000110","000110","010111","000110","000110","000110","010110","010110","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","010110","000110","101011","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","000110","000110","010110","010110","010101","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","000110","000110","000110","010110","010110","010110","010110","010101","010101","010101","010101","010100","010101","101001","011010","010110","000110","000110","000110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","010110","000110","000110","010110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010110","000110","000110","000110","010110","010110","000110","010110","010110","010101","010101","010101","010101","010101","010101","101001","101010","010101","000110","000110","000110","000110","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","000110","000110","000110","010110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","010111","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010110","000110","000110","000110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000110","000111","000110","010110","010101","101010","101110","010101","010101","010110","010110","000110","000110","000110","000110","000110","000110","000111","000110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010110","000110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","000110","000110","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010101","010101","010110","010101","010101","010101","010101","010101","010101","101001","111110","111001","111101","111101","111101","111101","111101","111110","010110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","000110","000110","000110","000110","000110","010110","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111001","010101","010110","010110","010101","010101","010101","010101","010101","101001","101010","111110","111101","111101","111101","111101","111101","111110","010101","010110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111001","101001","101001","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111001","010101","000110","000110","000110","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","010110","010110","010110","010101","010110","010110","000110","000110","000111","000110","000110","000110","000110","000110","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","010101","000110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","100100","011000","101001","111101","111101","111101","111101","111101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","010110","010110","000110","000110","000110","010110","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","100100","101001","101001","111101","111101","111101","111101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111101","010100","010110","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","010110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010101","010101","010101","010101","010101","010101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010101","011001","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111001","011001","010110","000110","000110","010110","010110","101111","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","010101","111110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","010110","010110","000111","000111","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","100100","010110","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000111","010110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","000111","000110","000110","000110","000110","010110","010110","010110","010110","010110","010101","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010101","000110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010110","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","011001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111001","010101","010110","000110","000110","010111","000110","000110","010101","010100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","000110","000110","000111","000111","000110","000110","010110","010101","010101","010101","010101","101000","111001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","010110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010110","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","000110","000110","000111","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","010110","010101","010101","101010","111101","111101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","010110","000110","000110","000110","010110","000000","101111","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011011","000110","000110","010110","010101","111110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010110","000111","000111","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","010110","000111","000110","000111","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","010110","000110","000111","010110","010110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010101","010110","000110","000110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","010110","000110","010110","010101","111110","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010110","000111","000111","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","000110","000110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011011","010110","000110","000110","010110","010110","010101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","010110","010110","010110","000110","010110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","010110","000110","000110","010101","101010","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111110","010110","000110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","000110","000110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","010110","000110","000110","000110","010110","000110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","000110","000110","000110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","111101","111101","101001","101001","010110","000110","000110","010110","010110","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","111101","111101","111001","101001","011001","010110","000110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010101","000110","000110","000110","000110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","010110","000110","010110","010110","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","010101","000110","000110","000111","000110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","010110","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","111101","111101","111101","101001","101001","010101","010101","010101","010101","010101","010110","000110","000111","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","111101","111101","111110","101001","011001","010101","010101","010101","010101","010101","010101","010110","000110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010101","010110","000110","000111","000111","000110","000110","010101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","010110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","010110","000110","000110","000110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","101010","010101","010110","010110","010110","000110","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","111101","101001","010101","010100","010101","010101","010101","010110","010110","010110","010110","010110","000110","000110","010110","000110","000110","010110","000110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111101","111101","101001","100100","010100","010101","010101","010101","010101","010110","010110","010110","000110","010110","000110","010110","000110","000110","000110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000111","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010101","010110","010110","010110","010110","010101","011001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010110","000110","000110","000110","101011","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111001","101001","010101","010101","010110","010110","000110","000110","000110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","011001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010100","010101","010101","010110","010110","010110","010110","010110","010110","010110","000110","000110","000110","000110","000110","010110","010110","010110","000110","000110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","010101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010100","010101","010101","010101","010110","010110","010110","010110","010110","010110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","011001","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","010110","010110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101000","010101","010101","010101","010101","101000","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","000110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","000110","010110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","011001","010101","010110","010110","010110","010110","000110","000110","000110","010110","000110","010110","101111","000000","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010110","000110","010110","010110","010110","101011","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010110","010101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","000110","000110","000110","010110","010110","011010","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","011001","010110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","111101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","011001","010101","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","000110","000110","010110","010101","111110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010101","010110","000110","000110","000110","000110","000110","000110","000110","000110","010110","101111","101111","101111","101011","010110","010110","010110","010110","010110","010110","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000111","000110","000110","000110","010110","010110","010110","010110","010110","010110","101011","101011","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","010101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010101","010110","010110","000110","000110","010110","010110","010110","010110","010110","010110","010110","011010","101011","101111","000000","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","011001","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","000110","010110","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111001","010101","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","000110","010110","010110","000110","010110","000110","000110","000110","000110","000110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","011010","101011","101111","000000","000000","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","010110","000110","000110","000110","011010","101111","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","011001","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","000110","000111","010110","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010101","000110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","101000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","000110","010111","000111","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","000110","000110","000110","000110","000110","010110","011010","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","010110","000110","101111","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011011","010110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","011001","010110","000110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","011001","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","010110","000110","000110","000111","000111","000111","000111","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010101","010110","010110","000110","000110","010110","010110","101111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010101","111001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","000110","011011","101011","101011","101011","101011","101011","101011","101011","101011","101011","101011","101011","101011","101011","101011","101011","101011","101011","101011","101011","101011","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010110","000110","000110","010111","000110","101011","101011","101111","101011","101011","101011","101011","101011","101011","101011","101011","101011","101011","101011","101011","101011","101011","101011","101011","101011","101011","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","000110","000101","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","000110","000110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010101","010110","000110","000110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010101","010101","010101","010101","010101","101001","101010","101110","010110","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010111","000110","000110","010110","000110","000110","000110","010110","010110","000110","010110","010110","000110","000110","000110","000110","010110","000110","000110","010110","010110","010110","000110","000110","000110","011010","000000","000000","000000","000000","000000","000000","000000","101111","000110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010110","000110","000111","000110","000110","000110","010110","000110","010110","000110","000110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","000110","010110","010110","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","010110","010110","010110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","000110","000110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","000110","000110","010101","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010101","010110","010110","010110","010101","010101","010101","010101","010101","010101","010100","010100","100100","101001","111001","111101","111101","111101","111101","111101","111101","111101","101010","010110","000110","000110","000110","010110","101111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010100","010101","000110","000110","000110","010110","000110","000110","010110","000110","000110","010110","000110","010110","010110","010110","010110","000110","000110","000110","010110","010110","010110","010110","010110","010110","000110","000110","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","010110","010110","010110","010110","000110","010110","010110","000110","010110","000110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","000110","010110","010110","000110","000110","010110","010110","000110","010110","101011","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","010110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","010110","000110","000110","010110","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","010110","010101","111110","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","101000","010100","010101","010101","011001","101001","111110","111110","111101","111101","111101","111101","111101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","000110","010101","101000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010100","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010110","000110","000110","000110","010110","010110","101111","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010110","000110","000110","010110","010110","010110","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","000110","010110","000110","000110","010110","011001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","010110","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111101","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","000110","010110","101011","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","000110","010101","101000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111001","101001","101001","111110","101010","111010","111110","101101","111001","111001","111001","101001","101001","101010","111010","101001","101001","101001","101001","101001","101010","111010","111001","101110","101110","101110","010110","000110","010110","000110","010110","101111","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111001","101101","101101","111010","101001","111010","101001","111010","101001","101001","111110","101010","101010","111110","101010","101010","101001","101101","101001","101010","101010","101110","101101","101001","101010","101010","011010","010110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","000110","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","010101","010110","010110","000110","000110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010110","000110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","000110","010101","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","010101","010110","000110","000110","010110","101011","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","010110","010110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010110","000110","000111","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","000110","000110","010110","010101","111110","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111001","010101","010110","010110","000110","000110","010110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","101011","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010101","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010110","000111","000111","000110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","010110","010101","010101","101001","111101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","010101","010101","010110","000110","000110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","010110","000110","000110","010110","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111110","010101","000110","000110","010110","010110","101010","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","101011","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010101","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011011","010110","000110","010110","000110","000110","010110","010101","010101","101001","111110","111110","111101","111101","111101","111101","111101","111101","111101","101001","010101","010101","010110","010110","010110","000110","000110","010110","011010","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","010110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","111101","111101","111101","101010","101010","010110","000110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","010110","000110","000110","010101","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010101","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","111110","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","101010","010101","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000110","000110","000110","010110","000110","000110","010110","010110","010101","010101","010101","010101","010101","010101","010101","010101","010101","010110","010110","000110","000110","000110","000110","000110","000110","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","111101","111101","111101","111101","101001","101001","010100","010100","010101","010101","010101","010110","010110","000110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","000110","000110","000110","010110","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","010101","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","010110","000110","000110","000110","000110","010110","010110","010101","010101","010101","010101","010101","010110","010101","010110","010110","010110","010110","000110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","010110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010110","010110","010110","000110","000110","000110","000110","000110","010110","010110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","010110","000110","000110","010110","010100","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","111101","111101","111101","111101","111110","101001","010101","010101","010101","010101","010101","010101","010110","010110","010110","010110","000110","000110","000110","000110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","010110","000110","000110","010110","101111","000000","000000","000000","000000","000000","010110","000110","000110","000110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010101","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","011010","010110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000111","000110","000110","000110","010110","010110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","000110","000110","000110","000110","000110","000110","010110","000110","000110","000110","000110","000110","000110","000110","000110","010110","000110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","010110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111101","111101","111101","111101","111101","111101","111101","101001","101001","010101","010101","010101","010101","010101","010101","010110","010110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","000110","010110","101111","000000","000000","000000","000000","000000","010110","000110","000110","010110","010101","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010110","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","101111","000110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","000110","000110","000110","000110","000110","010110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","010110","010110","000110","010110","010110","000110","010110","000110","010110","010110","010110","000110","010110","101010","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","010110","000110","000110","010110","010101","111110","111110","111101","111101","111110","101001","011001","010101","010101","010101","010101","010101","010110","010110","010110","010110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010110","010110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010101","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","000110","010110","101111","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","101111","000000","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","101111","101011","101011","101011","011010","101011","101011","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","010110","000110","000110","000110","000101","010101","010101","010101","010101","010101","010110","010110","010110","010110","000110","000110","000110","000110","000110","000111","000110","000110","000110","000110","000110","000110","010110","010110","000110","000110","000110","010110","010110","010110","010110","101011","101111","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010101","111110","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","010101","000110","000110","000110","010110","101111","000000","000000","000000","000000","000000","010110","000110","000110","000110","010110","101001","111101","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111101","101001","010110","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","000110","010110","000110","010110","010110","010110","000110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010110","010110","010110","011010","101011","101111","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","010110","010101","101110","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","101110","010110","000110","000110","010110","010110","101111","000000","000000","000000","000000","000000","010110","010110","000110","000110","010110","010101","111110","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111101","111110","010101","000110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","010110","000110","000110","000110","010110","000110","000110","000110","010110","010110","010110","000110","010110","010110","010110","000110","010110","010110","011011","101011","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","010110","000110","000110","010110","010110","010101","010110","010110","010110","010110","010101","010101","010101","010110","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010110","010110","010110","000110","000110","000110","010110","010110","000000","000000","000000","000000","000000","000000","101011","010110","000110","000110","000110","000110","010110","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010110","010110","010101","010101","010101","010101","010101","010101","010101","010101","010101","010101","010110","000110","000110","000110","000110","010110","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","000110","010110","010110","010110","000110","000110","010110","010110","010110","011011","101011","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011010","000110","010110","000110","000110","000110","000110","010110","000111","000111","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000111","000111","000110","000110","000110","010110","011010","000000","000000","000000","000000","000000","000000","000000","011010","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101011","011010","101011","101011","101111","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","010110","000110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","010110","000110","000110","000110","000110","000110","000110","000110","000110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","101011","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010110","000110","010110","000110","000110","010110","000110","010110","010110","000110","000110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","000110","010110","010110","010110","010110","010110","010110","010110","011010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","000000","000000","000000","000000","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"));


constant singleplayerString : singleplayer := (('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','1','1','1','1','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','0'),
('0','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1'),
('0','0','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','0','0','0'),
('0','0','0','1','1','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','1','0','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','1','1','1','1','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0'),
('0','1','1','1','0','0','0','1','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','0','0','0','0','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','0','0','0','1','1','1','0','0','0','0','0'),
('0','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0'),
('0','0','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));


constant multiplayerString : multiplayer :=(('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','1','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','1','1','1','1','1','1','1','1','1','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','0'),
('0','1','1','1','0','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','1','1','1','1','1','1','1','1','1','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1'),
('0','1','1','1','0','1','1','1','0','0','0','0','0','1','1','1','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','0','0','0'),
('0','1','1','1','0','1','1','1','1','0','0','0','0','1','1','1','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','1','0','0','0','0'),
('0','1','1','1','0','0','1','1','1','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','0'),
('0','1','1','1','0','0','1','1','1','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','0','0','0','0','0'),
('0','1','1','1','0','0','0','1','1','1','0','0','1','1','1','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','0','0','0','0','0'),
('0','1','1','1','0','0','0','1','1','1','0','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0'),
('0','1','1','1','0','0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0'),
('0','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0'),
('0','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','0','0','0','1','1','1','0','0','0','0','0'),
('0','1','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0'),
('0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','1','1','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','1','1','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));


constant NotString : Nott :=(('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0'),
('0','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0'),
('0','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0'),
('0','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','0'),
('0','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','0'),
('0','1','1','1','0','1','1','1','0','0','1','1','1','0','0','0','1','1','1','1','0','0','0','1','1','1','1','0','0','0','1','1','1','0','0','0','0'),
('0','1','1','1','0','0','1','1','1','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0'),
('0','1','1','1','0','0','1','1','1','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0'),
('0','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0'),
('0','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0'),
('0','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0'),
('0','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0'),
('0','1','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','0'),
('0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));


constant VeryEffectiveString : VeryEffective :=(('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0'),
('0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0'),
('0','0','1','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0'),
('0','0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0'),
('0','0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0'),
('0','0','0','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','1','1','0','1','1','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','0','1','1','1','1','1','1','1','1','0','0','1','1','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0'),
('0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0','0','0','0','0','1','1','1','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0'),
('0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','0','0','0','0','1','1','1','0','0','1','1','1','1','0','0','0','1','1','0','0','1','1','1','0','0','0','0','0','1','1','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0'),
('0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','0','0','0','1','1','1','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0'),
('0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','0','0','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','0','0','0','0','1','1','1','0','0','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0'),
('0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','0','0','0','0','0','0','1','1','1','0','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','0','0','0','0','1','1','1','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0'),
('0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','1','0','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','0','0','0','0','1','1','1','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0'),
('0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','0','0','1','1','1','0','0','0','0','1','1','0','0','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0'),
('0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','0','0','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0'),
('0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));


constant AustossFrontString : Pokemon :=(("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","111111","100110","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","100110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","100110","100110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","000000","111111","111111","100110","100110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","111111","111111","100110","100110","100110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","100110","100110","100110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","100110","100110","100110","100110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","010001","000000","000000","000000","000000","000000","010001","111111","111111","100110","100110","100110","111111","111111","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","100110","100110","100110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","111111","000000","010001","000000","000000","000000","000000","000000","000000","010001","111111","010001","100110","100110","100110","100110","010001","000000","000000","000000","000000","000000","111111","111111","111111","100110","100110","100110","100110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","010001","000000","000000","010001","010001","000000","000000","000000","000000","000000","111111","111111","100110","100110","100110","010001","100110","010001","100110","100110","100110","000000","100110","100110","100110","100110","100110","100110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","010001","000000","000000","000000","000000","000000","010001","010001","010001","000000","000000","000000","111111","010001","100110","100110","100110","010001","100110","100110","100110","100110","000000","010001","100110","100110","100110","100110","100110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","010001","100110","100110","010001","100110","010001","100110","000000","010001","010001","000000","010001","100110","100110","100110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","100110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100110","010001","100110","100110","100110","010001","100110","100110","111111","111111","100110","100110","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","010001","010001","010001","010001","000000","000000","000000","010001","100110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","010001","100110","100110","100110","100110","100110","100110","100110","100110","010001","010001","000000","100110","100110","100110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","100110","100110","010001","000000","000000","000000","000000","111111","010001","100110","100110","100110","100110","100110","100110","100110","100110","010001","010001","000000","010001","100110","010001","100110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","100110","100110","111111","111111","111111","111111","111111","000000","000000","000000","000000","010001","000000","000000","000000","100110","010001","010001","010001","000000","100110","111111","010001","100110","100110","100110","100110","100110","100110","100110","100110","010001","000000","100110","010001","100110","010001","000000","000000","100110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","100110","100110","100110","111111","111111","111111","111111","111111","111111","111111","111111","010001","000000","000000","100110","010001","010001","010001","000000","111111","010001","100110","100110","100110","100110","100110","100110","100110","100110","100110","100110","010001","100110","010001","100110","100110","100110","000000","100110","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100110","100110","100110","111111","111111","111111","100110","100110","100110","100110","010001","000000","010001","010001","010001","010001","000000","111111","111111","010001","100110","100110","100110","100110","100110","100110","100110","100110","100110","100110","100110","111111","111111","111111","000000","100110","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("010001","010001","010001","010001","010001","010001","010001","000000","000000","000000","000000","000000","000000","100110","100110","100110","100110","100110","100110","100110","100110","010001","000000","100110","010001","010001","010001","010001","000000","111111","111111","010001","010001","100110","100110","100110","100110","100110","010001","010001","010001","100110","100110","111111","111111","100110","000000","100110","000000","000000","000000","000000","000000","000000","000000","000000"),
("010001","100110","100110","111111","111111","111111","111111","111111","111111","000000","100110","000000","000000","000000","000000","100110","100110","100110","100110","100110","100110","010001","010001","100110","010001","010001","010001","010001","010001","000000","100110","111111","111111","010001","100110","100110","100110","100110","111111","111111","111111","010001","100110","100110","100110","100110","000000","100110","010001","000000","000000","000000","000000","000000","000000","000000"),
("000000","010001","000000","000000","100110","100110","100110","111111","111111","000000","100110","010001","000000","000000","000000","000000","000000","100110","100110","100110","010001","010001","010001","000000","111111","010001","010001","010001","010001","010001","000000","000000","100110","111111","111111","010001","100110","100110","100110","100110","111111","111111","010001","100110","100110","100110","000000","010001","100110","010001","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","100110","100110","100110","000000","100110","000000","000000","000000","000000","100110","000000","000000","010001","010001","010001","000000","000000","000000","111111","111111","100110","010001","010001","010001","010001","000000","000000","111111","111111","010001","100110","100110","100110","100110","100110","000000","100110","100110","010001","100110","000000","000000","100110","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","100110","000000","100110","000000","000000","000000","000000","100110","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","100110","100110","010001","010001","010001","010001","000000","111111","111111","010001","100110","100110","100110","100110","000000","100110","010001","100110","010001","010001","000000","010001","100110","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100110","000000","000000","000000","100110","010001","010001","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100110","100110","010001","010001","010001","000000","111111","010001","100110","100110","100110","000000","100110","010001","100110","010001","000000","010001","000000","100110","010001","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100110","010001","000000","000000","000000","100110","010001","010001","010001","000000","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","100110","100110","010001","010001","000000","100110","111111","010001","100110","100110","010001","100110","100110","010001","100110","000000","000000","000000","010001","100110","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","100110","010001","000000","000000","000000","000000","100110","010001","010001","000000","010001","100110","100110","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","100110","010001","010001","010001","000000","111111","010001","100110","100110","100110","100110","100110","100110","100110","111111","111111","000000","000000","010001","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","100110","010001","000000","000000","000000","000000","000000","100110","010001","000000","010001","100110","111111","111111","100110","010001","000000","000000","000000","000000","000000","100110","000000","000000","000000","100110","010001","010001","000000","100110","111111","100110","100110","111111","100110","111111","100110","100110","100110","111111","111111","111111","000000","000000","000000","010001","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","100110","010001","000000","000000","000000","000000","100110","010001","010001","000000","010001","100110","111111","111111","100110","010001","000000","000000","000000","100110","111111","111111","000000","000000","000000","100110","010001","010001","010001","000000","111111","010001","100110","100110","111111","100110","100110","100110","100110","100110","100110","111111","111111","111111","111111","100110","010001","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","010001","000000","000000","000000","000000","111111","010001","010001","000000","000000","000000","010001","100110","100110","010001","000000","000000","000000","100110","111111","111111","111111","000000","000000","000000","000000","100110","010001","010001","000000","111111","010001","100110","111111","100110","111111","100110","100110","100110","100110","100110","100110","100110","100110","100110","100110","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","010001","000000","000000","000000","000000","100110","010001","010001","000000","000000","000000","000000","010001","010001","000000","000000","000000","100110","111111","111111","111111","111111","000000","000000","000000","000000","100110","010001","010001","000000","111111","010001","100110","100110","111111","100110","111111","100110","100110","100110","100110","100110","100110","100110","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","100110","010001","000000","000000","000000","100110","010001","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","100110","111111","111111","111111","111111","111111","000000","000000","000000","000000","100110","010001","010001","000000","111111","010001","100110","100110","100110","111111","100110","100110","100110","100110","100110","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","100110","010001","000000","000000","000000","111111","010001","010001","010001","000000","111111","000000","000000","000000","000000","000000","100110","111111","000000","111111","111111","111111","000000","000000","000000","000000","000000","100110","010001","010001","100110","111111","100110","100110","100110","100110","100110","100110","100110","100110","010001","000000","010001","010001","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","100110","010001","000000","000000","000000","111111","010001","010001","010001","000000","111111","111111","100110","000000","000000","000000","000000","111111","000000","111111","111111","111111","000000","100110","100110","000000","000000","100110","010001","000000","111111","010001","100110","100110","100110","100110","010001","100110","100110","100110","010001","000000","010001","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","100110","010001","000000","000000","000000","100110","010001","010001","010001","000000","010001","111111","000000","000000","000000","000000","000000","000000","111111","111111","111111","000000","000000","111111","100110","000000","100110","010001","010001","100110","111111","010001","100110","100110","100110","100110","111111","010001","100110","010001","010001","000000","010001","010001","100110","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","100110","000000","000000","000000","000000","100110","010001","010001","000000","000000","100110","010001","000000","000000","000000","000000","000000","000000","000000","000000","010001","111111","111111","100110","000000","100110","010001","010001","111111","010001","100110","100110","100110","100110","100110","111111","111111","010001","010001","010001","000000","010001","010001","010001","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","100110","010001","000000","000000","000000","100110","010001","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100110","010001","111111","111111","000000","000000","100110","010001","000000","111111","010001","100110","100110","100110","100110","100110","100110","111111","000000","010001","010001","100110","000000","010001","010001","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","000000","100110","000000","000000","000000","000000","100110","010001","010001","000000","000000","000000","000000","000000","000000","000000","100110","010001","111111","111111","010001","111111","000000","000000","000000","100110","010001","100110","111111","100110","100110","100110","100110","100110","100110","100110","100110","000000","010001","100110","100110","000000","010001","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","010001","111111","100110","000000","100110","010001","000000","000000","000000","100110","010001","010001","010001","000000","000000","100110","111111","111111","111111","111111","010001","111111","100110","010001","000000","000000","000000","100110","010001","010001","111111","010001","100110","100110","100110","100110","100110","100110","000000","000000","100110","100110","000000","100110","000000","010001","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","100110","100110","100110","100110","000000","100110","010001","000000","000000","000000","100110","100110","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100110","010001","010001","111111","010001","100110","100110","100110","100110","100110","000000","010001","100110","100110","100110","111111","000000","000000","010001","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","100110","100110","000000","000000","000000","000000","100110","010001","000000","000000","000000","000000","100110","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","010001","010001","010001","100110","111111","010001","100110","100110","100110","100110","010001","100110","100110","100110","100110","111111","111111","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","000000","000000","000000","000000","100110","100110","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","010001","010001","010001","000000","111111","010001","100110","100110","100110","100110","100110","100110","100110","100110","100110","100110","111111","111111","111111","000000","010001","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100110","000000","000000","000000","000000","000000","000000","100110","010001","010001","010001","010001","000000","000000","000000","000000","000000","000000","100110","010001","010001","010001","000000","100110","111111","100110","100110","100110","100110","100110","100110","100110","100110","100110","100110","100110","100110","111111","111111","010001","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100110","010001","000000","000000","000000","000000","000000","100110","010001","010001","010001","010001","010001","010001","010001","010001","010001","010001","100110","010001","010001","010001","010001","000000","111111","010001","100110","100110","100110","100110","100110","010001","100110","100110","100110","100110","100110","100110","111111","111111","111111","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100110","010001","000000","000000","000000","000000","000000","000000","111111","010001","010001","010001","010001","010001","010001","010001","010001","010001","000000","100110","010001","010001","010001","000000","111111","010001","100110","100110","100110","100110","100110","100110","010001","010001","000000","000000","000000","100110","100110","111111","111111","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100110","010001","000000","000000","000000","000000","000000","000000","111111","100110","100110","100110","010001","010001","010001","010001","010001","010001","000000","100110","010001","010001","000000","111111","010001","100110","100110","100110","100110","100110","100110","010001","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100110","100110","010001","000000","000000","000000","000000","000000","000000","000000","000000","100110","100110","100110","010001","010001","010001","010001","010001","010001","000000","000000","111111","010001","100110","100110","100110","100110","100110","010001","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100110","100110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100110","010001","100110","100110","100110","010001","100110","010001","100110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100110","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100110","111111","010001","100110","100110","010001","100110","010001","100110","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","100110","100110","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","010001","100110","100110","100110","100110","010001","100110","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","100110","100110","100110","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","100110","100110","100110","100110","010001","100110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","100110","000000","000000","000000","000000","000000","000000","010001","000000","000000","000000","000000","000000","000000","010001","000000","000000","000000","000000","010001","010001","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","100110","000000","000000","000000","100110","010001","010001","010001","000000","010001","010001","010001","010001","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","100110","000000","000000","000000","000000","000000","100110","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"));

constant BisaflorFrontString : Pokemon :=(("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110001","111111","111111","110001","110001","110001","110001","110001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110001","110001","110001","110001","110001","110001","110001","111111","111111","110001","110001","110001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110001","110001","111111","111111","000000","000000","000000","000000","110001","110001","110001","110001","110001","110001","110001","110001","110001","110001","110001","110001","000000","000000","000000","000000","110001","110001","110001","110001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","110001","110001","110001","110001","110001","110001","110001","110001","110001","000000","110001","110001","000000","111111","000000","000000","111111","000000","110001","110001","000000","110001","110001","110001","110001","110001","110001","110001","110001","110001","110001","110001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110001","110001","110001","111111","111111","110001","110001","110001","110001","110001","110001","110001","110001","110001","000000","000000","111111","111111","111111","111111","111111","111111","000000","000000","110001","110001","110001","110001","111111","111111","110001","110001","110001","110001","110001","110001","110001","110001","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110001","110001","110001","110001","110001","110001","110001","110001","111111","111111","110001","110001","110001","110001","000000","111111","111111","000000","000000","000000","000000","111111","111111","000000","110001","110001","110001","110001","110001","111111","111111","110001","110001","110001","111111","111111","110001","110001","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","110001","000000","000000","110001","110001","110001","110001","110001","110001","111111","110001","110001","110001","000000","000000","110001","000000","000000","111111","111111","111111","111111","000000","000000","110001","000000","000000","110001","110001","110001","110001","110001","110001","110001","110001","110001","111111","111111","110001","110001","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110001","110001","110001","110001","110001","110001","110001","110001","000000","000000","000000","000000","110001","000000","000000","111111","000000","000000","111111","111111","000000","000000","111111","000000","000000","110001","110001","000000","000000","000000","110001","110001","110001","110001","110001","110001","110001","110001","110001","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","110001","110001","110001","110001","110001","110001","000000","000000","000000","110001","110001","110001","110001","110001","110001","110001","000000","000000","111111","111111","111111","111111","000000","000000","110001","110001","110001","110001","110001","110001","110001","000000","000000","000000","110001","110001","110001","110001","110001","110001","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110001","110001","110001","000000","000000","110001","110001","110001","110001","110001","110001","110001","110001","110001","110001","110001","110001","000000","000000","000000","000000","110001","110001","110001","111111","111111","110001","110001","110001","110001","110001","110001","110001","000000","000000","110001","110001","110001","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110001","000000","000000","110001","110001","110001","111111","111111","110001","110001","110001","110001","110001","111111","110001","110001","110001","110001","000000","110001","110001","110001","110001","110001","111111","110001","110001","110001","110001","110001","110001","110001","110001","110001","110001","000000","110001","110001","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110001","110001","110001","111111","111111","111111","111111","110001","110001","110001","111111","111111","110001","110001","110001","000000","000000","000000","000000","110001","110001","110001","110001","110001","110001","110001","110001","111111","111111","111111","110001","110001","110001","110001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110001","110001","110001","110001","111111","111111","110001","110001","110001","110001","110001","110001","110001","110001","110001","000000","000000","000000","000000","000000","000000","110001","110001","110001","110001","110001","110001","110001","110001","111111","111111","111111","110001","110001","110001","110001","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110001","110001","110001","110001","110001","110001","110001","110001","110001","110001","110001","110001","110001","110001","000000","000000","011101","011101","011101","011101","011101","011101","000000","110001","110001","110001","110001","110001","110001","110001","110001","110001","110001","110001","110001","110001","110001","110001","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110001","110001","110001","110001","110001","000000","110001","110001","110001","110001","110001","110001","000000","000000","000000","000000","111111","111111","011101","011101","000000","000000","000000","000000","110001","110001","110001","110001","110001","110001","000000","110001","110001","110001","110001","110001","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110001","110001","000000","110001","110001","110001","110001","110001","110001","000000","000000","011101","111111","111111","000000","000000","000000","000000","011101","011101","011101","000000","000000","110001","110001","110001","110001","110001","110001","000000","110001","110001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110001","110001","110001","110001","110001","110001","000000","000000","011101","111111","111111","111111","111111","111111","111111","011101","011101","011101","000000","000000","110001","110001","110001","110001","110001","110001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011101","011101","011101","011101","011101","000000","000000","110001","110001","110001","110001","000000","011101","000000","000000","000000","000000","111111","111111","111111","111111","011101","000000","000000","000000","011101","000000","110001","110001","110001","110001","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","011101","011101","000000","011101","011101","111111","111111","000000","000000","011101","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","000000","111111","111111","011101","011101","011101","000000","000000","011101","011101","000000","000000","000000","011101","000000","011101","011101","011101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","011101","011101","111111","000000","000000","011101","011101","011101","011101","011101","011101","000000","000000","011101","011101","111111","111111","000000","000000","000000","000000","000000","000000","000000","011101","000000","000000","000000","000000","000000","011101","011101","011101","011101","011101","011101","011101","000000","011101","011101","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","011101","011101","111111","000000","000000","011101","011101","011101","011101","011101","000000","011101","000000","000000","011101","011101","011101","111111","000000","000000","011101","011101","011101","011101","011101","011101","011101","000000","000000","000000","000000","011101","011101","011101","111111","111111","000000","000000","011101","011101","011101","011101","000000","000000","011101","011101","000000","000000","000000","000000","000000"),
("000000","000000","000000","011101","011101","011101","000000","011101","011101","011101","011101","011101","000000","011101","011101","000000","000000","011101","011101","011101","111111","000000","000000","011101","011101","011101","011101","000000","011101","011101","011101","000000","000000","000000","011101","011101","011101","011101","011101","011101","011101","011101","011101","111111","000000","000000","011101","011101","011101","011101","000000","000000","000000","000000","000000","000000"),
("000000","000000","011101","011101","011101","011101","011101","011101","011101","000000","011101","011101","000000","011101","000000","000000","000000","000000","011101","111111","000000","011101","011101","011101","011101","011101","011101","011101","000000","000000","011101","011101","000000","011101","011101","011101","000000","011101","011101","011101","011101","011101","011101","011101","011101","011101","111111","000000","000000","011101","011101","011101","011101","011101","000000","000000"),
("000000","000000","000000","011101","011101","000000","011101","011101","000000","011101","011101","000000","000000","000000","011101","011101","011101","011101","011101","000000","011101","011101","011101","011101","011101","000000","011101","011101","011101","011101","000000","000000","000000","000000","011101","000000","011101","011101","011101","000000","011101","011101","000000","011101","011101","011101","011101","011101","011101","000000","011101","011101","000000","011101","000000","000000"),
("000000","000000","000000","000000","000000","000000","011101","011101","000000","011101","011101","000000","000000","000000","011101","000000","011101","011101","000000","011101","011101","011101","000000","011101","011101","011101","000000","000000","011101","011101","000000","000000","000000","000000","000000","000000","000000","011101","000000","000000","011101","011101","000000","011101","011101","011101","000000","011101","011101","011101","011101","011101","011101","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011101","000000","011101","011101","011101","011101","011101","011101","011101","000000","011101","011101","011101","011101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011101","011101","000000","000000","011101","011101","000000","011101","011101","000000","011101","011101","011101","011101","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","111111","011101","011101","011101","000000","000000","011101","011101","011101","011101","011101","011101","011101","011101","011101","000000","011101","011101","000000","000000","000000","011101","011101","011101","000000","000000","000000","000000","000000","011101","011101","000000","011101","011101","000000","000000","011101","011101","000000","000000","011101","011101","000000","011101","011101","011101","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","110001","111111","111111","011101","011101","000000","011101","011101","000000","011101","011101","011101","000000","011101","011101","011101","000000","000000","000000","000000","011101","111111","111111","011101","000000","011101","000000","000000","011101","011101","011101","011101","011101","000000","000000","011101","000000","011101","011101","000000","000000","011101","011101","000000","000000","011101","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","110001","111111","111111","111111","000000","011101","011101","000000","011101","011101","011101","000000","000000","011101","011101","011101","000000","000000","000000","011101","111111","111111","011101","000000","110001","011101","000000","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","000000","000000","011101","000000","000000","000000","000000","011101","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","000000","011101","000000","000000","011101","011101","011101","000000","000000","011101","011101","011101","000000","011101","011101","011101","011101","011101","000000","110001","110001","011101","000000","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","000000","000000","000000","011101","011101","011101","000000","000000","000000","011101","011101","000000","000000","011101","011101","011101","011101","011101","011101","000000","000000","011101","011101","000000","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","000000","011101","011101","011101","011101","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","111111","111111","011101","111111","111111","111111","111111","000000","011101","011101","011101","000000","011101","000000","000000","000000","011101","011101","011101","000000","000000","011101","011101","011101","011101","011101","011101","011101","000000","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","111111","111111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","111111","011101","011101","111111","111111","111111","111111","000000","011101","011101","000000","011101","011101","011101","011101","011101","011101","011101","000000","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","000000","011101","011101","011101","011101","011101","011101","000000","011101","011101","011101","011101","011101","011101","000000","011101","111111","111111","011101","000000","000000"),
("000000","000000","000000","000000","000000","111111","000000","011101","011101","111111","111111","111111","111111","011101","000000","000000","000000","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","000000","011101","011101","011101","011101","011101","000000","011101","011101","011101","011101","011101","011101","011101","000000","011101","011101","011101","011101","011101","000000","011101","011101","111111","011101","000000","000000"),
("000000","000000","000000","000000","000000","111111","110001","000000","011101","111111","111111","111111","111111","111111","011101","011101","011101","011101","011101","011101","011101","011101","011101","000000","111111","111111","011101","000000","000000","000000","011101","011101","011101","011101","011101","011101","000000","011101","011101","000000","011101","011101","011101","011101","000000","011101","011101","011101","000000","011101","011101","011101","011101","011101","000000","000000"),
("000000","000000","000000","000000","111111","111111","110001","000000","011101","111111","111111","111111","111111","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","111111","000000","000000","110001","111111","000000","011101","011101","011101","011101","011101","011101","000000","011101","011101","011101","000000","011101","011101","011101","000000","011101","011101","011101","000000","011101","011101","011101","011101","011101","000000","000000"),
("000000","000000","000000","000000","111111","111111","111111","000000","111111","111111","111111","111111","111111","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","000000","000000","111111","000000","110001","111111","000000","011101","011101","011101","011101","011101","011101","011101","000000","011101","000000","011101","011101","011101","011101","011101","000000","011101","000000","011101","011101","011101","011101","011101","011101","000000","000000"),
("000000","000000","000000","011101","000000","111111","000000","111111","111111","111111","111111","111111","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","000000","111111","111111","111111","111111","011101","011101","011101","000000","011101","011101","011101","011101","000000","011101","011101","011101","011101","011101","011101","011101","000000","000000","011101","011101","011101","011101","011101","011101","000000","000000","000000"),
("000000","000000","000000","011101","000000","111111","111111","111111","111111","111111","111111","111111","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","000000","000000","011101","011101","011101","011101","000000","011101","011101","011101","011101","000000","011101","011101","011101","011101","011101","011101","011101","000000","000000","011101","011101","011101","011101","011101","000000","000000","000000","000000"),
("000000","000000","011101","111111","011101","000000","011101","111111","111111","111111","111111","111111","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","000000","011101","011101","011101","011101","000000","011101","011101","011101","011101","011101","000000","011101","011101","000000","011101","111111","000000","011101","111111","011101","011101","111111","000000","000000"),
("000000","000000","111111","111111","111111","000000","000000","011101","011101","111111","000000","111111","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","000000","000000","000000","011101","011101","011101","011101","011101","000000","011101","011101","011101","011101","011101","011101","000000","011101","011101","000000","000000","000000","111111","111111","011101","000000","000000","000000","000000"),
("000000","000000","111111","111111","111111","011101","000000","000000","000000","011101","011101","011101","011101","011101","000000","011101","011101","011101","011101","011101","011101","011101","011101","011101","000000","000000","000000","111111","110001","110001","000000","011101","011101","011101","000000","000000","011101","011101","011101","011101","011101","011101","000000","011101","011101","011101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","111111","111111","011101","011101","011101","011101","000000","000000","000000","011101","011101","011101","011101","011101","011101","011101","000000","000000","000000","000000","000000","110001","110001","110001","110001","110001","000000","011101","011101","011101","000000","000000","000000","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","011101","011101","011101","011101","011101","011101","000000","011101","000000","000000","000000","000000","000000","000000","110001","110001","110001","110001","110001","110001","110001","111111","000000","000000","011101","011101","011101","000000","000000","000000","000000","000000","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","111111","011101","011101","011101","011101","011101","011101","000000","000000","011101","011101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011101","011101","011101","011101","000000","000000","000000","000000","000000","000000","000000","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","011101","011101","011101","011101","011101","011101","000000","000000","000000","000000","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011101","011101","011101","011101","011101","011101","011101","011101","011101","011101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","111111","000000","011101","000000","111111","011101","000000","011101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011101","011101","011101","011101","011101","011101","011101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","011101","011101","111111","011101","011101","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"));

constant GallopaFrontString : Pokemon :=(("000000","000000","000000","000000","000000","000000","000000","000000","110000","110000","000000","110000","000000","000000","000000","000000","000000","000000","000000","110000","110000","000000","000000","000000","000000","110000","111100","110000","111100","000000","000000","000000","000000","111100","000000","000000","000000","111100","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111100","110000","110000","110000","110000","000000","000000","000000","000000","110000","110000","111100","111100","110000","110000","111100","110000","111100","110000","000000","000000","000000","111100","110000","111100","000000","000000","000000","111100","110000","111100","110000","000000","000000","000000","000000","111100","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","110000","111100","110000","110000","000000","000000","000000","110000","111100","111100","111100","111100","111100","111100","110000","110000","110000","111100","111100","111100","110000","110000","000000","000000","000000","000000","111100","110000","111100","110000","111100","110000","000000","000000","111100","110000","111111","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","110000","000000","000000","110000","111100","111100","110000","000000","000000","110000","111100","111100","111100","111100","111100","110000","110000","110000","110000","111100","111100","110000","110000","111100","000000","000000","000000","000000","000000","110000","111100","110000","111100","110000","110000","110000","111100","110000","110000","110000","000000","110000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","110000","000000","000000","110000","111100","111100","110000","110000","110000","000000","110000","111100","111100","110000","111100","110000","110000","110000","110000","110000","110000","110000","110000","110000","110000","000000","000000","000000","000000","000000","110000","111100","111100","110000","110000","110000","110000","110000","110000","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","110000","111100","110000","000000","110000","111100","110000","111100","110000","110000","110000","111100","111100","110000","111100","110000","111100","110000","110000","110000","110000","110000","110000","110000","000000","111100","110000","110000","110000","000000","110000","111100","111100","110000","110000","111100","110000","110000","110000","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","111100","111100","111100","110000","111100","111100","111100","110000","110000","111100","110000","111100","110000","111100","110000","110000","110000","110000","110000","111100","110000","111100","110000","110000","110000","110000","111100","110000","111100","111100","111100","111100","110000","110000","111100","000000","111100","110000","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","111100","110000","111100","111100","110000","111100","111100","110000","110000","110000","110000","111100","110000","110000","110000","110000","110000","111100","110000","111100","110000","111100","110000","111100","000000","110000","110000","110000","111100","111100","111100","111100","110000","111100","110000","000000","000000","000000","000000","000000","000000","000000","110000","110000","110000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","110000","111100","111100","110000","111100","111100","111100","110000","110000","110000","111100","110000","110000","110000","110000","110000","111100","110000","111100","110000","111100","111100","111100","111100","111100","000000","110000","110000","110000","111100","111100","111100","111100","110000","110000","110000","111100","000000","000000","000000","110000","111100","111100","111100","111100","110000","110000","110000","000000","000000","000000","000000","000000"),
("000000","000000","000000","110000","111100","111100","110000","111100","111100","111100","110000","110000","110000","110000","110000","110000","110000","110000","111100","110000","111100","110000","111100","110000","111100","111100","111100","111100","111100","111100","110000","111100","110000","111100","110000","110000","110000","110000","110000","111100","000000","110000","110000","111100","111100","111100","111100","111100","111100","111100","111100","110000","000000","000000","000000","000000"),
("000000","000000","000000","110000","111100","110000","111100","111100","111100","110000","111100","110000","110000","110000","110000","000000","000000","110000","110000","110000","110000","111100","110000","111100","110000","111100","110000","111100","111100","111100","111100","110000","111100","110000","110000","110000","000000","110000","111100","000000","110000","111100","111100","111100","111100","111100","110000","111100","110000","111100","110000","111100","110000","000000","000000","000000"),
("000000","000000","000000","000000","111100","110000","111100","111100","111100","111100","110000","110000","110000","110000","000000","111100","111100","110000","110000","110000","110000","110000","110000","110000","110000","110000","111100","110000","111100","111100","110000","111100","110000","110000","110000","000000","000000","000000","000000","000000","110000","111100","111100","111100","111100","110000","111100","110000","111100","110000","111100","110000","110000","000000","000000","000000"),
("000000","000000","000000","000000","110000","110000","111100","110000","111100","110000","110000","110000","110000","000000","111100","110000","111100","000000","110000","110000","110000","110000","110000","110000","110000","110000","110000","111100","111100","110000","111100","110000","111100","110000","110000","000000","000000","000000","000000","000000","110000","111100","111100","111100","110000","111100","110000","110000","110000","110000","110000","110000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","110000","111100","110000","111100","110000","110000","000000","111100","110000","110000","111100","000000","110000","110000","110000","110000","110000","110000","110000","110000","110000","110000","110000","111100","110000","110000","110000","110000","111100","000000","000000","000000","000000","000000","000000","110000","111100","110000","111100","110000","110000","110000","110000","111100","110000","110000","110000","000000","000000","000000"),
("000000","110000","000000","000000","000000","000000","000000","110000","111100","110000","110000","110000","000000","111100","110000","110000","111100","000000","110000","110000","000000","110000","000000","110000","110000","110000","110000","110000","110000","110000","110000","111100","110000","111100","110000","000000","000000","000000","000000","000000","000000","110000","110000","110000","110000","110000","110000","110000","111100","110000","111100","110000","111100","110000","110000","000000"),
("110000","111111","111111","111111","000000","000000","111111","000000","110000","110000","110000","000000","111100","110000","110000","110000","111100","000000","110000","110000","110000","000000","110000","000000","110000","110000","110000","110000","110000","110000","110000","111100","110000","110000","110000","110000","111100","111111","000000","000000","110000","110000","110000","110000","110000","110000","111100","111100","110000","111100","110000","111100","110000","111100","110000","110000"),
("000000","000000","111100","111100","111111","111111","111100","110000","110000","000000","000000","111100","111100","110000","110000","111100","000000","110000","000000","000000","000000","000000","110000","110000","110000","110000","110000","110000","110000","110000","111100","110000","110000","110000","111100","111111","111111","111111","111111","111111","000000","110000","110000","000000","110000","110000","110000","111100","111100","110000","110000","110000","110000","110000","111100","110000"),
("000000","000000","000000","111100","111100","111100","000000","000000","000000","111111","111111","111100","111100","111100","111100","000000","111100","111100","111100","111111","111111","111100","111100","000000","000000","110000","110000","110000","110000","111100","110000","110000","111100","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","110000","111100","111100","110000","110000","110000","110000","110000","111100","110000","110000"),
("000000","110000","000000","000000","000000","000000","111111","111111","111100","111100","111100","111111","111100","111100","111100","111100","111100","111100","111100","111100","111100","111111","111111","111100","111111","111100","000000","000000","111100","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111100","000000","000000","000000","000000","110000","110000","110000","110000","110000","110000","110000","110000","000000"),
("110000","111111","111111","111100","111100","111100","111100","111100","111100","111100","111111","111100","111111","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111111","111100","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111100","111111","111100","000000","000000","000000","110000","110000","110000","110000","111100","111100","110000","000000","000000"),
("000000","110000","000000","000000","111100","111100","111100","111100","111100","111100","111100","111111","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111111","111100","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111100","111111","000000","000000","000000","000000","110000","110000","111100","111100","110000","110000","000000","000000"),
("000000","000000","000000","000000","110000","000000","000000","111100","111100","111100","111111","111111","111111","111100","110000","000000","111100","111100","110000","111100","111100","111100","111100","111100","111100","111111","111100","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111100","111111","111100","000000","000000","000000","000000","110000","111100","111100","110000","110000","000000","000000","000000"),
("000000","000000","000000","000000","000000","111111","111111","110000","111100","111111","111111","111111","111111","110000","000000","111100","111100","111100","000000","111100","111100","111100","111100","111100","111100","111100","111111","111100","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111100","111111","111100","110000","000000","110000","111100","111100","111100","110000","110000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111100","000000","110000","111111","111100","111100","111100","110000","111100","111100","111100","111100","111100","111100","111100","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111100","111100","000000","000000","110000","111100","111100","111100","110000","110000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111100","000000","110000","000000","111100","111100","111100","000000","111100","111100","111100","111100","111100","111100","111111","111100","111111","111111","111111","111111","111111","111111","111111","111111","111100","111111","111111","111111","111111","111111","111100","111100","111100","000000","000000","110000","111100","111100","111100","111100","110000","110000","000000","000000"),
("000000","000000","000000","000000","000000","110000","111100","111111","111111","111111","111111","111111","111100","111100","000000","111100","111100","111100","111100","000000","111100","111100","111100","111100","111100","111100","111100","111111","111111","111111","111111","111111","111111","111111","111111","111100","110000","111111","111111","111111","111111","111111","111100","111100","111100","000000","000000","000000","110000","111100","110000","111100","111100","110000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111100","111100","111100","111100","111100","111100","000000","111100","111100","111100","111100","111100","111100","111111","111100","111111","111111","111111","111111","111111","111111","111111","111111","000000","111111","111111","111111","111111","111111","111100","111100","111100","110000","000000","000000","110000","111100","110000","110000","110000","111100","110000","000000"),
("000000","000000","000000","000000","000000","000000","110000","111100","111111","111111","111111","111111","111111","111100","111100","111100","111100","111100","111100","110000","111100","111100","111100","111100","111100","111100","111100","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","111111","111111","111111","111111","111111","111100","111100","000000","000000","000000","000000","000000","110000","110000","110000","110000","110000","110000","110000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111100","111100","111100","111100","111100","000000","111100","111100","111100","111100","111100","111100","111100","111111","111100","111111","111111","111111","111111","111111","111111","111111","111111","000000","111100","111111","111111","111111","111100","111100","111100","000000","000000","000000","000000","000000","000000","000000","110000","110000","110000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111100","111100","111100","111100","111100","000000","111111","111100","111100","111100","111100","111100","111100","111111","111100","111111","111111","111111","111111","111111","111111","111111","111111","111100","000000","000000","111111","111111","111111","111100","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111100","111100","111100","111100","111100","000000","110000","111111","111100","111100","111100","111100","111111","111100","111111","111111","111111","111111","111111","111111","111111","111100","111100","111100","000000","000000","111100","111111","111111","111100","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","110000","110000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111100","111100","111100","111100","000000","110000","111100","110000","000000","111100","111100","111100","111100","111111","111100","111111","111111","111111","111111","111111","111100","111100","111100","000000","000000","000000","000000","111111","111100","111111","111100","111100","000000","000000","110000","110000","000000","000000","110000","110000","110000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","110000","111111","111111","111111","111100","111100","000000","111100","111100","000000","111100","110000","111100","110000","111100","111100","111100","111111","111100","111111","111111","111111","111111","111111","111111","111100","111100","000000","000000","000000","000000","000000","111100","111111","111100","111100","111100","000000","000000","111100","110000","110000","110000","111100","110000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","110000","111111","111100","111111","111100","000000","111100","111100","000000","110000","000000","000000","110000","111100","110000","111100","111100","111100","111111","111111","111111","111111","111111","111111","111111","000000","111100","000000","000000","000000","000000","000000","000000","111100","111111","111100","111100","111100","000000","110000","111100","110000","111100","110000","111100","110000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111100","111100","111100","111100","000000","000000","110000","111100","110000","000000","110000","110000","110000","110000","111111","111100","111111","111111","111111","111111","111111","111111","111100","000000","000000","000000","000000","000000","000000","000000","000000","111100","111100","111100","110000","110000","111100","110000","110000","110000","110000","110000","110000","110000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110000","111100","110000","111100","110000","000000","000000","110000","110000","110000","110000","111100","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","110000","110000","111100","111100","111100","110000","110000","110000","110000","110000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110000","111111","111111","111111","000000","111100","110000","111100","110000","111100","000000","110000","000000","000000","110000","000000","111100","111111","111111","111111","111111","111111","111111","000000","000000","000000","111100","000000","000000","000000","000000","000000","111100","111100","110000","110000","111100","110000","110000","110000","110000","110000","110000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","110000","111111","111111","000000","111111","111100","111100","111100","111100","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111100","000000","000000","000000","000000","111100","000000","000000","000000","000000","111100","111100","111100","111100","110000","110000","000000","000000","110000","110000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","110000","111111","111100","000000","111111","111111","111100","111100","111100","110000","000000","000000","000000","000000","000000","000000","000000","111100","111111","111111","111111","111111","111100","000000","000000","110000","000000","110000","111100","000000","000000","000000","000000","111100","111100","110000","110000","110000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111100","110000","111111","111111","110000","000000","111111","111100","111100","111100","110000","000000","000000","000000","000000","000000","000000","000000","000000","111100","111111","111111","111111","111111","000000","111100","110000","111100","110000","111100","000000","000000","000000","000000","000000","111100","111100","110000","110000","110000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","110000","110000","111100","110000","000000","111111","111111","111100","111100","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","000000","110000","111100","110000","111100","111100","110000","000000","000000","000000","000000","111100","111111","110000","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","110000","111100","110000","000000","111111","111111","111111","111100","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","111111","111111","111100","110000","111100","111100","111100","111100","110000","110000","000000","000000","000000","000000","111111","110000","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111100","110000","110000","000000","111111","111111","111111","111100","000000","110000","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","111111","111111","110000","111100","111100","111100","111100","110000","111100","110000","000000","000000","000000","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","110000","110000","000000","111111","111111","111100","111100","000000","000000","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110000","111111","111111","111100","111100","110000","111100","110000","111100","110000","111100","000000","000000","110000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","110000","110000","000000","111100","111100","111100","110000","111100","000000","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111100","111100","110000","110000","110000","110000","110000","111100","000000","000000","000000","000000","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","110000","110000","000000","111100","111100","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","111111","110000","110000","110000","110000","110000","110000","000000","000000","000000","000000","000000","111111","000000","000000","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","110000","000000","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111100","111100","110000","110000","110000","110000","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110000","111111","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","111100","110000","110000","110000","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110000","000000","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110000","111111","111100","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111100","111100","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110000","110000","111100","111100","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110000","000000","000000","000000","000000","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"));

constant GaradosFrontString : Pokemon :=(("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","000000","111111","111111","111111","111111","000000","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111100","000000","111111","111111","111111","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111100","000000","111111","000000","111111","111111","111100","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","111100","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111100","000000","000000","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","000000","111111","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111100","000000","000000","111111","111100","111100","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111100","111111","000000","111111","111100","000000","000000","010111","010111","111111","000000","000000","111111","111111","111111","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","111111","111100","111111","111100","111100","000000","010111","010111","111111","111111","111111","111111","000000","000000","111111","111111","111100","000000","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111100","111111","111100","111111","000000","010111","010111","111111","010111","111111","111111","000000","000000","000000","000000","000000","000000","000000","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111100","000000","010111","010111","010111","111111","010111","010111","010111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","111111","111111","111111","111111","111111","111100","000000","010111","010111","010111","010111","010111","010111","111111","010111","111111","111111","111111","111111","111111","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","010111","000000","111111","111111","111111","111100","000000","010111","010111","010111","010111","010111","010111","111111","010111","111111","111111","111111","111111","010111","010111","010111","000000","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","111111","010111","000000","000000","000000","000000","000000","000000","000000","010111","010111","000000","000000","010111","111111","010111","111111","111111","111111","010111","010111","010111","000000","000000","010111","010111","010111","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","111111","111111","111111","111111","010111","111111","010111","010111","000000","000000","000000","010111","000000","010111","010111","111111","111111","010111","010111","010111","000000","000000","010111","010111","010111","010111","010111","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","000000","111111","111111","111111","111111","010111","010111","010111","010111","000000","010111","000000","000000","010111","010111","010111","010111","010111","000000","000000","000000","010111","010111","010111","010111","010111","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","111111","111111","111111","111111","010111","010111","010111","000000","010111","000000","000000","010111","010111","010111","010111","010111","000000","010111","010111","000000","010111","010111","010111","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","000000","111111","111111","010111","010111","010111","000000","010111","010111","000000","010111","000000","010111","010111","010111","000000","010111","010111","000000","010111","010111","010111","010111","000000","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","000000","010111","010111","010111","000000","000000","010111","010111","000000","000000","010111","000000","010111","010111","010111","010111","010111","010111","000000","010111","010111","010111","000000","111100","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","010111","000000","010111","010111","000000","000000","010111","000000","010111","000000","010111","000000","000000","010111","010111","010111","000000","010111","010111","010111","000000","000000","000000","000000","000000","010111","000000","010111","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","010111","010111","000000","010111","000000","000000","000000","010111","000000","010111","000000","000000","010111","010111","010111","010111","010111","000000","000000","111111","111111","111111","111111","010111","010111","000000","010111","010111","010111","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","000000","010111","000000","000000","000000"),
("000000","010111","010111","000000","000000","000000","000000","000000","000000","000000","010111","000000","000000","000000","000000","010111","000000","000000","000000","010111","010111","010111","010111","010111","111111","111111","111111","111111","111111","010111","010111","010111","000000","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","111111","111100","000000","010111","000000","000000","000000"),
("111111","000000","000000","010111","010111","010111","000000","000000","000000","000000","010111","010111","000000","000000","010111","000000","000000","000000","111111","000000","010111","010111","010111","010111","111111","111111","111111","010111","010111","010111","010111","000000","000000","000000","010111","010111","010111","010111","010111","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","111111","111100","000000","010111","000000","000000","000000"),
("111111","111111","111111","000000","000000","000000","010111","010111","000000","000000","000000","010111","000000","000000","000000","000000","000000","111111","111111","111111","000000","010111","010111","111111","010111","111111","010111","010111","010111","000000","000000","000000","010111","010111","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","111100","111100","000000","010111","000000","000000","000000","000000"),
("111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","010111","010111","000000","000000","000000","111111","000000","111111","111111","000000","010111","010111","010111","111111","010111","010111","000000","000000","000000","010111","010111","010111","000000","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","111100","000000","010111","111100","111100","000000","010111","000000","000000","000000","000000"),
("111111","111111","111111","111111","111111","000000","010111","000000","010111","111111","000000","010111","010111","000000","000000","000000","000000","000000","010111","010111","010111","010111","010111","010111","010111","010111","000000","010111","000000","010111","010111","000000","000000","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","111111","000000","010111","010111","111100","000000","010111","000000","000000","000000","000000","000000"),
("111111","111111","111111","000000","000000","111111","010111","010111","000000","111111","111111","000000","010111","000000","000000","010111","010111","010111","000000","010111","010111","010111","010111","010111","010111","010111","010111","000000","010111","010111","000000","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","010111","111100","111111","000000","010111","010111","000000","010111","010111","000000","000000","000000","000000","000000"),
("111111","111111","000000","111111","111111","010111","010111","010111","000000","111111","000000","111111","000000","000000","010111","010111","000000","010111","010111","000000","010111","010111","010111","010111","000000","010111","000000","010111","010111","000000","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","010111","111100","111100","000000","111111","010111","010111","010111","000000","000000","000000","000000","000000","000000"),
("111111","111111","000000","010111","010111","010111","000000","010111","010111","000000","010111","010111","010111","010111","010111","000000","010111","000000","000000","000000","000000","010111","010111","010111","000000","000000","010111","010111","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","111111","010111","000000","000000","000000","010111","000000","000000","000000","000000","000000","000000","000000","000000"),
("111111","111111","111111","000000","000000","010111","010111","000000","010111","000000","010111","000000","000000","010111","010111","000000","000000","111100","111100","111100","111100","000000","010111","010111","000000","000000","010111","010111","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","111111","010111","010111","000000","000000","010111","010111","000000","000000","000000","000000","000000","000000"),
("111111","000000","000000","000000","000000","000000","000000","000000","010111","010111","010111","010111","000000","000000","000000","111100","111100","111100","000000","000000","111100","111100","000000","010111","010111","000000","010111","000000","111111","111111","111111","111111","010111","010111","010111","010111","010111","010111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","010111","010111","010111","010111","010111","000000","000000","000000","010111","000000","000000","111111","111111","111100","111100","111100","000000","111111","111111","000000","111100","111100","000000","010111","000000","010111","000000","111111","010111","010111","010111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","111100","111100","111100","000000","010111","000000","000000","000000","000000","000000"),
("000000","000000","111111","111111","000000","000000","010111","010111","000000","111100","111100","111100","111100","111100","111100","000000","000000","000000","010111","111111","000000","000000","111100","000000","010111","010111","000000","000000","010111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","000000","010111","000000","000000","000000","000000"),
("000000","000000","000000","111111","111111","111111","111111","000000","000000","000000","111100","010111","000000","000000","000000","000000","000000","000000","000000","010111","000000","000000","000000","111100","000000","010111","000000","111111","111111","111111","111111","111111","111111","111111","000000","000000","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","111100","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","111111","111111","111111","111111","111111","111111","000000","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","000000","000000","000000","111111","111111","111111","111111","111111","111111","000000","010111","010111","010111","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","000000","000000","111111","111111","000000","010111","000000","000000","000000"),
("000000","000000","000000","000000","111111","111111","111111","111111","111111","010111","000000","000000","111111","000000","000000","000000","000000","000000","000000","000000","010111","010111","000000","111100","000000","111111","000000","000000","111111","111111","111111","111111","111111","111111","000000","010111","010111","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","000000","111111","000000","000000","010111","111100","000000","000000","000000"),
("000000","000000","000000","000000","111111","111111","111111","010111","010111","111111","111111","000000","000000","111100","000000","000000","000000","000000","010111","010111","010111","010111","010111","000000","111100","000000","111111","111111","000000","111111","111111","111111","111111","111111","111111","000000","010111","010111","000000","000000","000000","000000","111111","010111","000000","000000","000000","000000","000000","000000","010111","010111","010111","010111","000000","000000"),
("000000","000000","000000","000000","111111","010111","010111","111111","111111","111111","111111","111111","000000","111100","000000","000000","000000","010111","010111","010111","010111","010111","010111","000000","111100","000000","000000","000000","111111","000000","111111","111111","000000","000000","000000","010111","010111","010111","000000","000000","000000","111111","111111","010111","111111","000000","000000","000000","000000","000000","010111","010111","000000","000000","000000","000000"),
("000000","000000","000000","000000","010111","111111","111111","111111","111111","111111","111111","000000","111111","000000","000000","000000","010111","010111","010111","010111","010111","010111","010111","010111","111100","000000","111100","111100","000000","111111","000000","000000","111100","111100","010111","010111","010111","010111","000000","000000","000000","111111","111111","010111","111111","000000","000000","000000","000000","000000","000000","000000","010111","010111","111100","010111"),
("000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","010111","111111","000000","111100","000000","010111","010111","010111","010111","010111","010111","010111","010111","000000","111100","000000","111100","000000","111111","000000","111100","111100","111100","111100","010111","010111","010111","000000","000000","111100","111111","111111","111111","111100","000000","000000","000000","000000","000000","000000","010111","010111","010111","111100","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","111111","000000","000000","111100","000000","010111","010111","010111","010111","010111","010111","010111","010111","000000","111100","000000","111100","000000","111111","000000","111100","111100","111100","111100","010111","010111","000000","010111","000000","111100","111111","111111","111111","000000","111111","000000","000000","000000","000000","000000","000000","000000","010111","010111","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","111111","000000","000000","000000","111100","010111","010111","010111","010111","010111","010111","010111","010111","000000","111100","000000","111100","000000","111111","000000","111100","111100","111100","010111","000000","000000","111100","111100","010111","000000","111111","111111","111111","111100","111100","000000","000000","000000","010111","000000","010111","010111","000000","010111","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","111111","000000","000000","000000","111100","000000","010111","010111","010111","010111","010111","000000","000000","000000","111100","000000","111111","111100","000000","111111","000000","111100","000000","000000","010111","000000","111100","111100","010111","000000","111111","111111","111100","111111","000000","000000","000000","000000","000000","010111","010111","010111","010111","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","111111","000000","000000","000000","000000","111100","000000","000000","000000","010111","010111","000000","111111","000000","000000","111100","000000","111100","111111","000000","111111","000000","000000","111100","010111","000000","111111","000000","010111","010111","010111","000000","111100","111111","111100","000000","000000","000000","000000","000000","010111","010111","010111","111100","010111","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","111111","000000","000000","000000","000000","111111","111111","000000","000000","000000","000000","000000","111111","000000","111100","111100","000000","000000","000000","000000","111111","000000","111100","111100","111100","000000","111111","000000","010111","010111","010111","000000","000000","111100","000000","000000","000000","000000","010111","010111","000000","000000","111100","111100","010111","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","010111","111111","010111","000000","000000","000000","000000","000000","111100","111100","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","111111","000000","010111","010111","010111","010111","000000","010111","111100","000000","000000","000000","010111","010111","010111","010111","010111","000000","010111","010111","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","111100","010111","000000","000000","000000","111100","111100","111100","111100","010111","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","000000","111100","010111","010111","010111","010111","000000","010111","000000","000000","010111","010111","000000","010111","010111","111100","010111","010111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","000000","000000","111100","111100","111100","111100","111100","000000","000000","010111","000000","000000","000000","010111","000000","000000","111100","000000","000000","000000","000000","111100","111100","010111","010111","010111","000000","111100","111100","010111","000000","111100","111100","010111","000000","111100","111100","111100","010111","010111","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","000000","000000","010111","000000","000000","000000","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","111111","111100","111100","111100","111100","010111","010111","000000","111100","111100","111100","000000","111100","111100","111100","010111","000000","111100","010111","010111","010111","000000","000000"),
("000000","000000","000000","000000","111111","000000","000000","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","111100","000000","000000","000000","111100","111100","111100","111100","111100","010111","000000","010111","010111","111100","010111","000000","111100","111100","010111","010111","000000","010111","010111","010111","000000","000000","000000"),
("000000","000000","000000","000000","000000","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","111111","111100","111100","111100","010111","000000","010111","010111","010111","010111","010111","000000","010111","010111","010111","010111","010111","000000","010111","010111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111100","111100","111100","000000","000000","010111","010111","010111","010111","010111","010111","000000","010111","010111","010111","010111","010111","000000","010111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","000000","000000","000000","111111","111100","111100","010111","010111","010111","010111","000000","010111","010111","010111","010111","010111","010111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","111111","111111","111111","111100","111111","111100","111100","111100","010111","010111","000000","010111","010111","010111","010111","010111","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","111111","111111","111100","111111","111100","111100","111100","000000","111100","111100","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","111111","111111","111111","000000","000000","111100","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"));

constant GlurakFrontString : Pokemon :=(("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","110100","000000","000000","000000","000000","111111","111111","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000000","000000","000000","000000","000000","000000","111111","111111","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111111","111111","111111","110100","110100","000000","000000","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","000000","000000","000000","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111111","000000","110100","000000","111111","111111","111111","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","000000","000101","000101","000101","000000","000000","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","111111","111111","110100","110100","000000","000000","000000","110100","000000","000000","111111","000000","111111","111111","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","000000","000101","000101","000101","000101","000101","000000","110100","110100","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","111111","111111","110100","000000","110100","110100","110100","110100","110100","110100","000000","000101","000000","111111","111111","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","000000","000101","000101","000101","000101","000101","000101","000000","110100","110100","000000","000000","000000","000000","000000","000000"),
("000000","110100","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","000000","000101","000101","000101","000101","000101","000101","000101","000000","110100","110100","000000","000000","000000","000000","000000"),
("000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","000000","000101","000101","000101","000101","000101","000101","000101","000101","000000","110100","000000","000000","000000","000000","000000"),
("000000","000000","110100","110100","000000","111111","000000","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","000000","000000","000000","000000","000000","110100","000000","000101","000101","000101","000101","000101","000101","000101","000101","000000","110100","110100","000000","000000","000000","000000"),
("000000","000000","111111","000000","000000","111111","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","000000","000000","000000","000000","110100","000000","000101","000101","000101","000101","000101","000101","000101","000101","000101","000000","110100","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","110100","000101","000101","000000","000000","000000","000000","000000","110100","110100","110100","110100","000000","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","000000","000000","110100","110100","000000","000101","000101","000101","000101","000101","000101","000101","000101","000101","000000","110100","110100","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","110100","000101","000101","000000","000000","110100","110100","110100","000000","000000","110100","110100","000000","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","000000","110100","110100","110100","000000","110100","000000","000101","000101","000101","000101","000101","000101","000101","000101","000101","000101","000101","000000","110100","000000","000000","000000"),
("000000","000000","000000","000000","000000","110100","000101","000101","000101","000000","110100","110100","110100","000000","000000","110100","110100","110100","000000","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","000000","110100","110100","000000","000000","000000","000101","000101","000101","000101","000101","000101","000101","000101","000101","000000","110100","000000","000000","000000"),
("000000","000000","000000","000000","000000","110100","000101","000101","000000","110100","111111","110100","110100","000000","110100","110100","000000","000000","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","000000","110100","110100","000000","000101","000101","000000","000000","000000","000101","000101","000101","000101","000101","000101","000101","000000","110100","110100","000000","000000"),
("000000","000000","000000","000000","110100","000000","000000","000000","000000","111111","111111","110100","000000","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","000000","110100","000000","000101","000101","000101","000101","000101","000000","000000","000101","000101","000101","000101","000101","000101","000101","000000","110100","000000","000000"),
("000000","000000","000000","000000","110100","000000","111111","000000","110100","111111","110100","110100","000000","110100","110100","000000","000000","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","000000","000101","000101","000101","000101","000101","000101","000000","000000","000101","000101","000101","000101","000101","000101","000000","110100","000000","000000"),
("000000","000000","000000","000000","110100","000000","000000","000000","110100","110100","110100","000000","000000","110100","000000","000101","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","000000","000101","000101","000101","000101","000101","000101","000101","000101","000000","000101","000101","000101","000101","000101","000101","000000","110100","000000","000000"),
("000000","000000","000000","000000","110100","000101","000000","000000","000000","110100","000000","000000","110100","110100","000000","000101","000101","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","110100","110100","000000","000101","000000","000101","000101","000101","000101","000101","000101","000101","000101","000000","000101","000101","000101","000101","000101","000000","110100","110100","000000"),
("000000","000000","000000","110100","110100","000101","000000","000000","000000","000000","110100","110100","110100","000000","000101","000101","000101","000000","110100","111111","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","110100","110100","110100","110100","000000","000101","000000","000101","000000","000101","000101","000101","000101","000101","000101","000101","000101","000101","000101","000101","000101","000101","000101","000000","110100","000000"),
("000000","000000","000000","110100","000101","000101","000101","000000","110100","110100","110100","000000","000000","000101","000101","000101","000101","000000","110100","110100","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000101","000000","000101","000101","000101","000101","000101","000101","000101","000101","000000","000000","000000","000101","000101","000101","000101","000000","110100","000000"),
("000000","000000","000000","110100","000101","000101","000101","000101","000000","000000","000000","000101","000101","000101","000101","000101","000000","000101","000000","111111","110100","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000101","000000","000101","000000","000000","000000","000000","000000","000101","000101","000000","110100","110100","000000","000000","000101","000101","000101","000000","110100","000000"),
("000000","000000","000000","110100","000101","000101","000000","000000","000000","000000","000000","000000","000000","000000","000101","000000","000101","000000","000000","110100","111111","110100","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","111111","000000","000000","000000","110100","110100","000000","000000","000000","000101","000101","000000","110100","000000"),
("000000","000000","000000","110100","000101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000000","000101","000000","111111","110100","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","110100","110100","110100","110100","111111","111111","111111","110100","110100","110100","110100","000000","000000","000000","000000","000101","000000","110100","000000"),
("000000","000000","000000","110100","000101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000000","000101","000000","111111","110100","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","110100","110100","110100","110100","111111","111111","111111","110100","110100","110100","110100","000000","000000","000000","000000","000101","000000","110100","000000"),
("000000","000000","000000","110100","000000","000000","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000101","000000","000000","110100","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","110100","110100","110100","110100","111111","111111","111111","000000","000000","110100","000000","000000","000000","000000","000000","000000","110100","110100","000000"),
("000000","000000","000000","111111","000000","000000","000000","000000","000101","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","110100","110100","110100","110100","111111","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","110100","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","110100","110100","000000","000000","110100","110100","110100","110100","000000","000000","110100","110100","110100","000000","000000","000000","000000","000000","110100","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","110100","110100","000000","111111","111111","000000","000000","000000","000000","111111","111111","110100","000000","110100","111111","111111","111111","111111","000000","000000","110100","000000","000000","110100","110100","110100","110100","110100","000000","110100","110100","000000","000000","000000","110100","110100","110100","110100","000000","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","111111","000101","110100","110100","000000","111111","111111","000000","000000","000000","000000","110100","110100","110100","000000","111111","111111","111111","111111","000000","111111","111111","000000","110100","110100","000000","110100","110100","110100","110100","000000","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111111","110100","110100","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","000000","000000","110100","000000","000000","110100","110100","110100","110100","000000","111111","111111","111111","111111","000000","111111","110100","110100","110100","110100","000000","110100","110100","110100","110100","000000","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","111111","110100","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","000000","110100","110100","000000","000000","111111","111111","111111","111111","111111","000000","000000","110100","110100","110100","110100","000000","000000","110100","110100","000000","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","110100","111111","110100","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","000000","000000","000000","111111","111111","111111","111111","000000","111111","000000","110100","110100","110100","110100","110100","110100","110100","110100","000000","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","110100","111111","110100","110100","110100","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","000000","000000","000000","000000","111111","111111","111111","111111","000000","111111","111111","110100","110100","110100","110100","110100","110100","110100","110100","000000","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111111","110100","110100","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","000000","000000","000000","000101","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","110100","110100","110100","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","111111","110100","110100","110100","110100","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","110100","110100","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","111111","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","111111","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","110100","110100","111111","111111","111111","110100","110100","110100","110100","110100","110100","000000","000000","000000","110100","110100","110100","110100","110100","110100","110100","111111","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","110100","110100","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","110100","111111","111111","111111","111111","111111","110100","110100","110100","110100","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","111111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","110100","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","110100","110100","111111","111111","111111","111111","111111","110100","110100","110100","110100","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","111111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","110100","110100","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","110100","110100","110100","111111","111111","111111","110100","110100","110100","110100","110100","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","110100","110100","110100","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","110100","110100","110100","110100","110100","110100","111111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","110100","110100","110100","110100","110100","111111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","000000","111111","111111","111111","111111","110100","111111","110100","111111","110100","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","110100","110100","110100","110100","111111","111111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","000000","000000","111111","110100","111111","110100","111111","110100","111111","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","110100","110100","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","000000","000000","110100","111111","110100","111111","110100","111111","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","000000","000000","000000","110100","000000","110100","110100","110100","000000","000000","000000","110100","111111","110100","111111","000000","000000","110100","110100","110100","110100","110100","110100","000000","000000","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","000000","000000","000000","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","110100","000000","000000","110100","000000","000000","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","000000","111111","111111","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","110100","110100","111111","111111","000000","110100","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","000000","111111","111111","000000","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"));

constant KokoweiFrontString : Pokemon :=(("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","111111","111111","111111","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","111111","111111","111111","111111","111111","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","001000","111111","111111","111111","111111","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","001000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","111111","001000","111111","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","001000","001000","001000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","001000","001000","001000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","001000","001000","001000","000000","000000","000000","111111","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","001000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","000000","000000","001000","001000","001000","000000","000000","111111","111111","001000","001000","111111","001000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","000000","001000","001000","001000","000000","000000","111111","001000","111111","111111","001000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","000000","001000","001000","000000","000000","001000","001000","111111","111111","111111","000000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","000000","000000","000000","000000","001000","001000","001000","001000","001000","000000","001000","000000","001000","001000","001000","001000","111111","000000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","001000","001000","001000","001000","000000","001000","000000","001000","001000","001000","001000","000000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","001000","001000","001000","001000","000000","000000","001000","001000","001000","000000","001000","001000","001000","001000","001000","001000","000000","000000","000000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","001000","111111","111111","111111","111111","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","001000","001000","001000","000000","001000","001000","001000","000000","001000","001000","001000","001000","001000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","001000","001000","001000","111111","001000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","001000","001000","000000","001000","001000","000000","000000","001000","001000","001000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","000000","000000","000000","000000","001000","001000","000000","001000","001000","001000","000000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","000000","000000","000000","000000","000000","001000","000000","000000","111111","111111","111111","111111","000000","000000","001000","001000","001000","000000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","100100","000000","001000","000000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","100100","100100","000000","001000","001000","000000","000000","000000","000000","111111","111111","100100","100100","000000","000000","000000","000000","000000","000000","001000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","100100","000000","111111","000000","111111","111111","000000","111111","111111","111111","100100","100100","000000","001000","000000","000000","000000","111111","111111","111111","111111","111111","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","100100","100100","000000","001000","000000","001000","111111","111111","001000","000000","000000","000000","001000","100100","100100","000000","000000","000000","111111","111111","001000","001000","001000","111111","111111","100100","001000","001000","000000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","001000","000000","000000","000000","001000","000000","000000","000000","000000","111111","000000","000000","100100","100100","000000","111111","111111","111111","111111","111111","100100","111111","111111","111111","111111","100100","100100","000000","000000","000000","111111","001000","111111","000000","111111","111111","111111","100100","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","111111","111111","100100","000000","100100","111111","000000","111111","111111","111111","111111","100100","000000","111111","111111","100100","100100","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","100100","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","100100","100100","100100","100100","100100","000000","111111","111111","111111","111111","111111","111111","111111","100100","111111","100100","111111","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","111111","111111","111111","111111","111111","000000","111111","111111","100100","001000","000000","000000","000000","000000","001000","111111","111111","111111","111111","100100","100100","000000","111111","111111","111111","000000","111111","111111","000000","000000","000000","000000","000000","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","001000","111111","111111","000000","001000","000000","111111","000000","000000","000000","000000","111111","000000","000000","001000","111111","100100","100100","000000","111111","111111","111111","111111","000000","001000","111111","111111","111111","111111","111111","000000","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","100100","000000","111111","111111","000000","000000","000000","001000","001000","000000","000000","111111","111111","111111","100100","100100","000000","100100","111111","111111","111111","111111","111111","001000","001000","001000","001000","001000","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","100100","111111","100100","111111","000000","111111","111111","111111","111111","001000","001000","001000","000000","111111","111111","111111","111111","100100","100100","000000","100100","100100","111111","100100","111111","100100","111111","100100","111111","100100","111111","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","000000","100100","111111","100100","111111","100100","111111","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","100100","100100","000000","000000","000000","100100","100100","111111","100100","111111","100100","111111","100100","111111","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","100100","100100","111111","100100","111111","100100","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","100100","100100","000000","000000","000000","100100","111111","100100","111111","100100","111111","100100","111111","100100","111111","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","100100","111111","100100","111111","100100","000000","111111","111111","111111","111111","111111","111111","111111","111111","100100","100100","000000","001000","001000","001000","000000","100100","111111","100100","111111","100100","111111","100100","111111","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","100100","100100","100100","100100","100100","000000","100100","111111","111111","111111","111111","100100","100100","100100","000000","001000","001000","100100","100100","100100","000000","100100","100100","100100","100100","100100","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","100100","100100","100100","000000","000000","000000","000000","001000","100100","100100","100100","100100","000000","000000","001000","100100","100100","000000","000000","000000","000000","000000","000000","100100","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","100100","100100","100100","100100","100100","100100","100100","000000","000000","000000","000000","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","100100","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","000000","000000","100100","100100","100100","000000","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","000000","111111","111111","000000","100100","100100","000000","100100","100100","100100","000000","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","100100","100100","100100","100100","100100","100100","100100","000000","100100","100100","100100","000000","100100","100100","000000","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","000000","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","100100","100100","100100","100100","100100","100100","100100","100100","000000","100100","100100","100100","000000","100100","000000","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","100100","100100","100100","100100","111111","111111","111111","100100","100100","100100","100100","100100","100100","000000","100100","000000","100100","100100","100100","100100","100100","100100","100100","100100","100100","100100","000000","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","100100","111111","111111","111111","111111","111111","100100","100100","000000","100100","100100","000000","100100","000000","100100","100100","100100","100100","100100","100100","100100","100100","100100","000000","100100","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","111111","111111","111111","111111","111111","100100","100100","000000","100100","000000","100100","000000","100100","100100","100100","100100","100100","100100","100100","100100","000000","000000","100100","100100","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","111111","111111","111111","111111","111111","100100","100100","000000","100100","000000","000000","000000","000000","000000","100100","100100","100100","100100","000000","000000","100100","100100","100100","100100","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","111111","111111","111111","111111","111111","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","111111","111111","111111","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","100100","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","000000","100100","100100","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","100100","000000","000000","000000","000000","000000","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","100100","100100","100100","100100","100100","100100","100100","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100100","000000","100100","000000","100100","100100","100100","000000","100100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","000000","100100","000000","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"));

constant MagmarFrontString : Pokemon :=(("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","000000","000000","100000","100000","100000","100000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","100000","100000","000000","000000","000000","100000","111111","100000","100000","111111","111111","100000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","100000","000000","000000","100000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","100000","100000","100000","111111","111111","100000","000000","000000","100000","111111","111000","111111","111000","111111","100000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","100000","000000","000000","100000","100000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","111111","111000","111111","111000","111111","100000","000000","000000","100000","111000","111000","111000","111000","111111","111000","100000","100000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","100000","100000","100000","100000","100000","100000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","111111","111000","111111","100000","000000","000000","000000","100000","111000","111000","111000","111000","111000","111000","111000","100000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","111000","100000","100000","100000","100000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","100000","111000","111000","111000","100000","000000","000000","000000","000000","100000","111000","111000","111000","111000","111000","111000","100000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","100000","111000","100000","100000","100000","100000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","111000","111000","111000","111000","111000","111000","100000","000000","000000","000000","000000","111000","111000","111000","111000","100000","100000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","000000","111000","100000","100000","111000","111000","111000","100000","100000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","111000","111000","111000","111000","100000","000000","000000","000000","000000","111000","100000","000000","000000","000000","000000","000000","000000","000000","100000","100000","100000","100000","100000","100000","111000","111000","100000","100000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","111000","100000","000000","000000","100000","100000","100000","000000","000000","100000","111000","100000","111000","100000","100000","000000","000000","000000","000000","100000","100000","000000","000000","000000","000000","000000","000000","000000","000000","100000","100000","100000","111000","100000","100000","100000","100000","100000","100000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","111000","100000","111000","100000","100000","111000","111000","111000","100000","100000","100000","100000","111000","100000","111000","000000","000000","000000","000000","100000","100000","100000","000000","000000","000000","000000","000000","000000","000000","000000","100000","100000","100000","100000","100000","111000","100000","100000","100000","100000","100000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","100000","100000","000000","100000","111000","111111","111111","111111","111000","100000","100000","100000","100000","111000","100000","000000","000000","000000","000000","100000","100000","100000","000000","000000","000000","000000","111000","000000","000000","000000","100000","100000","100000","100000","111000","111000","111000","100000","100000","100000","100000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","111000","100000","000000","100000","111000","111111","111111","111111","111111","111111","111000","100000","100000","100000","100000","100000","000000","000000","000000","100000","100000","100000","100000","000000","000000","000000","111000","100000","000000","000000","000000","000000","100000","100000","111000","100000","111000","100000","111000","100000","100000","100000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","111111","111000","100000","000000","100000","111000","111111","111111","111111","111111","111000","111000","100000","100000","100000","100000","100000","100000","000000","100000","100000","100000","100000","100000","000000","000000","100000","100000","100000","000000","000000","000000","000000","100000","100000","100000","111000","100000","111000","100000","111000","100000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","111111","111111","111000","100000","100000","000000","100000","100000","111000","111000","111000","111000","100000","100000","100000","100000","100000","100000","100000","100000","000000","000000","100000","100000","000000","000000","000000","000000","100000","100000","100000","000000","000000","000000","000000","000000","100000","100000","100000","100000","100000","111000","100000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","111111","111111","111111","111000","100000","100000","000000","100000","100000","100000","100000","100000","100000","100000","100000","100000","100000","100000","100000","100000","100000","100000","100000","000000","000000","111000","111000","111000","111000","000000","000000","000000","000000","100000","000000","000000","000000","000000","000000","100000","100000","111000","100000","111000","100000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","111000","111000","111000","100000","100000","100000","100000","000000","100000","100000","100000","100000","100000","100000","100000","100000","100000","100000","100000","100000","100000","100000","000000","111000","111000","111111","111111","111111","111000","111000","111000","000000","100000","100000","000000","100000","000000","000000","000000","000000","000000","100000","111000","100000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","100000","100000","100000","100000","100000","100000","100000","000000","000000","000000","000000","100000","100000","100000","100000","100000","000000","100000","100000","100000","100000","100000","100000","000000","111111","111111","111111","111111","111111","111000","111000","000000","100000","100000","100000","100000","100000","000000","000000","000000","000000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","100000","100000","100000","100000","100000","000000","000000","111111","111111","111111","111111","000000","000000","000000","000000","100000","100000","100000","100000","100000","100000","000000","111000","111111","111111","111111","111111","111111","111000","111000","111000","000000","100000","000000","100000","100000","000000","100000","000000","000000","100000","111000","111000","111000","100000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","100000","100000","111111","000000","111000","111000","000000","111111","000000","111111","111111","000000","100000","100000","100000","100000","100000","100000","000000","000000","111000","111000","111000","111111","111111","111111","111000","111000","111000","111000","000000","000000","000000","100000","100000","000000","100000","000000","000000","000000","111000","111000","111000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","111111","111000","111000","000000","000000","000000","000000","100000","100000","100000","100000","100000","100000","000000","000000","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","100000","100000","100000","100000","100000","000000","000000","000000","000000","111000","111000","111000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111000","111000","111000","111000","100000","100000","100000","100000","100000","100000","100000","100000","000000","000000","000000","100000","000000","111000","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000","100000","000000","000000","100000","100000","100000","100000","000000","111000","111000","111000","111000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111000","111000","111000","111000","111000","111000","111000","111000","000000","100000","100000","100000","100000","000000","000000","000000","100000","000000","111000","111000","111000","111000","111000","111000","111000","111000","000000","111000","000000","000000","100000","100000","100000","100000","100000","100000","100000","000000","000000","111000","111000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111000","000000","000000","111111","111000","111000","111000","111000","111000","111000","111000","000000","100000","100000","100000","000000","000000","000000","100000","100000","100000","000000","000000","111000","111000","111000","111000","000000","000000","100000","111000","000000","100000","100000","100000","100000","100000","100000","100000","000000","111111","111111","000000","111000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111000","100000","000000","000000","111000","111000","111000","111000","111000","111000","000000","100000","100000","000000","000000","000000","000000","000000","100000","100000","100000","100000","100000","000000","000000","000000","000000","100000","111000","111000","111000","000000","000000","000000","100000","100000","100000","100000","000000","000000","111000","111000","111111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","100000","100000","000000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","100000","100000","100000","100000","100000","100000","100000","100000","100000","100000","100000","100000","111000","111000","000000","111000","111111","000000","000000","000000","100000","000000","111111","111000","000000","000000","000000","111000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","111000","000000","100000","100000","100000","100000","100000","100000","100000","100000","111000","111000","100000","100000","111000","111000","111000","111000","000000","111111","000000","000000","111000","111111","000000","000000","111111","111111","000000","111000","111000","111000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","100000","100000","100000","111000","100000","100000","100000","100000","111000","111000","111000","111000","111000","111000","000000","000000","000000","111000","000000","111000","111111","000000","000000","000000","111111","000000","111000","111000","111000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","100000","100000","100000","100000","111000","100000","100000","100000","111000","111000","111000","111000","111000","000000","111000","111000","111000","111000","111000","000000","111111","000000","111000","000000","000000","111000","111000","111000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","111000","100000","100000","100000","111000","111000","100000","100000","100000","111000","111000","111000","111000","000000","111000","111000","111111","111111","111111","111000","000000","111000","111000","111000","000000","111000","111000","111000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","111000","000000","111000","111000","100000","111000","111000","111000","100000","100000","111000","111000","111000","111000","000000","111000","111000","111111","111111","111111","111111","111111","111000","111000","111000","111000","111000","100000","111000","111000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","111000","111000","111000","111000","100000","100000","111000","111000","111000","111000","111000","111000","111000","111000","000000","111000","111000","111111","111111","111111","111111","111111","111000","111000","111000","111000","111000","000000","111000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","100000","000000","111000","111000","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","111000","111000","111111","111111","111111","111111","111111","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","100000","100000","100000","100000","000000","111000","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","111000","111000","111000","111111","111111","111111","111000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","100000","100000","100000","000000","111000","111000","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","100000","100000","100000","100000","000000","111000","111000","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","100000","100000","100000","000000","000000","000000","000000","111000","000000","100000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","111000","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","111000","111000","111000","111000","111000","111000","000000","000000","000000","000000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","100000","100000","100000","000000","000000","000000","100000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","100000","100000","100000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","000000","100000","100000","100000","100000","100000","100000","100000","100000","100000","100000","100000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","000000","000000","000000","100000","100000","100000","100000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","100000","000000","000000","100000","100000","100000","100000","100000","100000","100000","000000","000000","000000","000000","000000","000000","000000","000000","100000","100000","100000","100000","100000","100000","100000","100000","100000","100000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","111111","111000","111000","000000","000000","111111","111111","000000","100000","100000","100000","100000","100000","100000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100000","100000","100000","100000","100000","100000","000000","000000","100000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","000000","000000","111111","111111","111000","111000","000000","100000","100000","100000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","100000","100000","100000","100000","000000","111111","111000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111000","000000","100000","100000","100000","000000","111111","111111","111111","111000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111000","000000","000000","000000","000000","000000","000000","111111","111111","111000","100000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"));

constant SarzeniaFrontString : Pokemon :=(("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110101","000000","000000","000000","000000","000000","110101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","000000","000000","110101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","011100","011100","000000","000000","111111","111111","011100","000000","000000","000000","000000","000000","011100","111111","111111","111111","000000","110101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","011100","011100","011100","011100","000000","111111","111111","011100","000000","000000","011100","011100","011100","011100","011100","000000","000000","000000","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","011100","011100","011100","011100","011100","011100","000000","111111","011100","000000","000000","011100","011100","011100","011100","011100","011100","011100","011100","000000","111111","000000","000000","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","111111","011100","111111","011100","111111","011100","011100","011100","000000","111111","011100","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","111111","011100","111111","011100","111111","011100","111111","011100","011100","111111","011100","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","011100","111111","011100","111111","011100","111111","011100","111111","000000","111111","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","011100","111111","011100","111111","011100","111111","011100","111111","011100","000000","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","111111","111111","110101","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","011100","111111","011100","111111","011100","111111","011100","011100","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","011100","111111","011100","111111","011100","111111","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","111111","111111","111111","011100","011100","011100","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","011100","011100","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","110101","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","111111","011100","011100","011100","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110101","110101","110101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110101","000000","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110101","110101","110101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","110101","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110101","110101","000000","000000","011100","011100","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","000000","110101","110101","110101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110101","000000","111111","000000","011100","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","000000","000000","000000","110101","110101","110101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110101","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","000000","000000","110101","110101","110101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","110101","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110101","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","000000","110101","110101","110101","110101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110101","110101","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","110101","110101","110101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110101","110101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110101","110101","110101","000000","000000","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110101","110101","110101","110101","000000","000000","000000","000000","000000","000000","110101","110101","110101","110101","110101","110101","000000","000000","000000","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110101","110101","111111","111111","110101","110101","110101","110101","110101","110101","110101","110101","110101","000000","000000","000000","000000","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110101","110101","111111","111111","111111","111111","110101","110101","110101","110101","000000","000000","111111","000000","000000","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110101","110101","110101","110101","110101","110101","000000","000000","000000","111111","111111","000000","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","111111","000000","000000","000000","111111","111111","000000","111111","000000","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","011100","011100","011100","011100","000000","000000","000000","011100","011100","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","111111","011100","111111","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","110101","000000","000000","000000","000000","011100","011100","011100","011100","011100","000000","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","000000","000000","011100","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","011100","111111","011100","011100","011100","011100","011100","000000","000000","111111","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","011100","000000","000000","011100","011100","000000","000000","000000","011100","011100","011100","011100","011100","011100","011100","000000","011100","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","110101","000000","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","011100","011100","011100","011100","000000","000000","111111","111111","111111","111111","111111","111111","011100","011100","011100","111111","011100","000000","011100","011100","011100","011100","011100","011100","011100","000000","000000","011100","111111","011100","111111","011100","011100","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","111111","111111","011100","000000","000000","000000","111111","011100","011100","011100","011100","011100","000000","000000","000000","011100","011100","000000","111111","111111","111111","111111","111111","111111","111111","011100","011100","111111","011100","000000","011100","011100","011100","011100","011100","011100","011100","111111","011100","000000","011100","111111","011100","111111","011100","011100","000000","000000","000000","000000","000000","000000"),
("000000","000000","110101","111111","111111","000000","000000","111111","011100","111111","011100","111111","011100","011100","011100","011100","011100","011100","011100","000000","011100","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","011100","011100","011100","011100","011100","111111","011100","111111","011100","111111","011100","000000","011100","111111","011100","111111","011100","011100","000000","000000","000000","000000","000000"),
("000000","000000","000000","111111","000000","011100","111111","011100","111111","011100","111111","011100","011100","011100","011100","011100","011100","011100","011100","011100","000000","111111","111111","011100","011100","011100","111111","111111","111111","111111","111111","111111","000000","011100","011100","011100","011100","111111","011100","111111","011100","111111","011100","111111","011100","011100","011100","111111","011100","111111","011100","000000","000000","000000","000000","000000"),
("000000","000000","011100","011100","011100","011100","011100","111111","011100","111111","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","000000","111111","111111","011100","011100","011100","111111","111111","111111","111111","111111","111111","011100","000000","000000","011100","011100","011100","111111","111111","111111","011100","111111","011100","111111","011100","000000","011100","111111","011100","011100","011100","000000","000000","000000","000000"),
("000000","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","000000","111111","111111","011100","011100","111111","111111","111111","111111","111111","111111","111111","111111","011100","111111","000000","000000","011100","011100","111111","111111","111111","111111","111111","011100","111111","011100","000000","011100","111111","011100","011100","000000","000000","000000","000000"),
("000000","011100","011100","011100","000000","000000","000000","000000","000000","000000","011100","011100","011100","011100","011100","011100","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","011100","111111","011100","011100","011100","000000","011100","011100","111111","111111","111111","011100","111111","011100","111111","000000","111111","011100","011100","011100","000000","000000","000000","000000"),
("000000","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","011100","111111","011100","111111","011100","000000","000000","000000","011100","011100","111111","111111","111111","011100","111111","011100","011100","000000","011100","011100","011100","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","011100","011100","111111","111111","111111","011100","111111","011100","011100","000000","000000","000000","000000","011100","011100","111111","111111","111111","011100","111111","011100","000000","011100","011100","011100","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","011100","011100","011100","111111","111111","011100","111111","011100","111111","011100","000000","000000","000000","000000","000000","011100","011100","111111","011100","011100","011100","011100","000000","011100","011100","011100","011100","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110101","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","011100","011100","111111","111111","011100","111111","011100","111111","011100","000000","000000","000000","000000","000000","000000","000000","011100","011100","111111","011100","011100","011100","011100","000000","011100","011100","011100","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","000000","110101","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","011100","111111","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","011100","111111","011100","011100","011100","011100","000000","011100","011100","011100","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","000000","110101","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","011100","111111","011100","111111","011100","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","011100","011100","011100","011100","000000","011100","011100","011100","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","011100","111111","011100","111111","011100","111111","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","011100","011100","011100","000000","011100","011100","011100","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","111111","011100","111111","011100","111111","011100","111111","011100","111111","011100","111111","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","011100","011100","011100","011100","011100","011100","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","110101","011100","111111","111111","111111","111111","111111","111111","011100","000000","000000","000000","000000","111111","011100","111111","011100","111111","011100","111111","011100","111111","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","000000","011100","011100","011100","011100","011100","011100","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","111111","111111","111111","111111","111111","011100","000000","000000","000000","000000","000000","000000","011100","111111","011100","111111","011100","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","000000","000000","011100","011100","011100","011100","011100","011100","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110101","011100","011100","011100","111111","111111","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","000000","000000","000000","011100","011100","011100","011100","011100","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","000000","000000","000000","000000","011100","011100","011100","011100","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110101","011100","011100","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","000000","000000","000000","000000","000000","000000","011100","011100","011100","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","000000","000000","000000","000000","000000","000000","000000","011100","011100","011100","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110101","000000","000000","000000","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"));

constant TurtokFrontString : Pokemon :=(("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","010111","000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","000000","010111","000000","000000","000000","000000","111111","111111","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","111111","010111","000000","000000","111111","111111","111111","010111","000000","000000","111111","111111","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","000000","000000","000000","111111","111111","111111","000000","111111","000000","000000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","010111","111111","000000","000000","000000","000000","000000","111111","111111","111111","111111","000000","000000","000000","000000","000000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","010111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","111111","010111","010111","111111","111111","111111","111111","000000","000000","000000","000000","000000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","000000","111111","000000","000000","010111","010111","111111","010111","111111","010111","000000","000000","000000","000000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","000000","111111","111111","000000","010111","010111","111111","010111","111111","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","111111","111111","010111","000000","000000","010111","111111","010111","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","010111","000000","000000","000000","000000","000000","010111","000000","000000","111111","111000","111000","111000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","111111","111111","010111","010111","010111","010111","000000","000000","000000","010111","111111","111111","111111","111111","010111","000000","000000","111000","111111","000000","000000","010111","010111","111111","111111","000000","000000","000000","000000","000000","111111","111000","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","010111","010111","010111","010111","010111","010111","010111","000000","000000","000000","111111","111111","111111","111111","111111","111111","000000","000000","010111","111111","111111","111000","111111","111000","111111","111000","000000","000000","111111","111111","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","000000","000000","111111","111111","111111","111111","111111","111111","000000","111111","111000","111111","111000","111111","111000","111000","111111","111111","111111","111111","111111","010111","000000","000000","000000","010111","111000","111000","111000","111000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","010111","111111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","000000","000000","000000","000000","000000","000000","111111","000000","111111","111000","111111","111000","111000","000000","111111","111111","111111","010111","000000","000000","000000","000000","000000","000000","000000","010111","111000","111000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","010111","111111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","111111","111111","111111","111111","010111","010111","000000","111111","010111","111000","111000","111000","111000","000000","111111","111111","000000","000000","000000","010111","111111","111111","010111","010111","000000","000000","010111","111000","111000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","010111","111111","010111","111111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","111111","111111","111111","010111","000000","010111","000000","111111","000000","111000","111000","111000","111000","111000","000000","000000","000000","000000","111111","111111","000000","000000","000000","000000","010111","000000","000000","111000","111000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","111111","010111","111111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","000000","000000","010111","000000","111111","111111","010111","111000","111000","111000","111000","111000","010111","000000","111111","111111","000000","000000","000000","000000","000000","000000","010111","000000","010111","111000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","111111","010111","010111","010111","010111","010111","010111","111111","111111","111111","010111","010111","010111","010111","010111","010111","000000","000000","000000","010111","000000","111111","111111","000000","111000","111000","111000","111000","111000","000000","010111","111111","000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","111000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","010111","010111","010111","010111","010111","010111","111111","111111","111111","010111","010111","010111","010111","000000","010111","010111","010111","000000","000000","010111","000000","111111","111111","111111","010111","111000","111000","111000","010111","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","000000","010111","010111","010111","010111","010111","010111","111111","111111","111000","010111","010111","000000","000000","010111","010111","010111","010111","010111","010111","010111","000000","111111","111111","111111","000000","111000","111000","111000","000000","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","010111","010111","010111","010111","010111","000000","111000","010111","010111","000000","000000","111111","111111","000000","010111","010111","010111","010111","010111","010111","000000","010111","111111","111000","000000","111000","111000","010111","000000","000000","111111","111111","010111","000000","000000","000000","000000","000000","000000","000000","010111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","010111","010111","010111","010111","010111","010111","010111","010111","000000","000000","000000","111111","000000","111111","111111","000000","010111","010111","010111","010111","010111","010111","000000","000000","111000","111111","000000","111000","111000","000000","000000","000000","010111","111111","111111","000000","000000","000000","000000","000000","000000","010111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","010111","000000","111111","111111","000000","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","000000","000000","000000","111111","111111","010111","010111","010111","010111","010111","010111","000000","000000","000000","111111","111000","111111","000000","111000","000000","000000","000000","010111","111111","111111","111111","000000","000000","000000","000000","010111","010111","000000","000000","000000","000000"),
("000000","000000","000000","000000","111111","111111","111111","000000","111111","000000","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","000000","000000","000000","111000","111111","111000","000000","010111","000000","000000","010111","000000","010111","111111","111111","111111","111111","111111","111111","010111","000000","000000","000000","000000","000000"),
("000000","000000","000000","111111","111111","010111","010111","000000","010111","010111","010111","010111","010111","000000","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","000000","000000","000000","111111","111000","111111","000000","000000","000000","010111","000000","010111","000000","010111","010111","111111","111111","111111","010111","000000","111000","000000","000000","000000","000000"),
("000000","010111","111111","111111","010111","111111","010111","010111","000000","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","000000","010111","010111","010111","010111","000000","000000","000000","111000","111111","111000","010111","000000","000000","000000","010111","000000","010111","000000","000000","010111","010111","010111","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","111111","010111","111111","010111","010111","010111","010111","000000","000000","000000","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","000000","010111","010111","010111","000000","000000","000000","010111","111111","111000","111111","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","111000","000000","000000","000000","000000"),
("000000","111111","111111","111111","010111","111111","010111","010111","010111","010111","000000","111000","000000","000000","000000","000000","000000","000000","000000","010111","010111","010111","010111","010111","010111","000000","111000","111000","010111","000000","000000","000000","000000","111111","111000","111111","111000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","111000","000000","000000","000000","000000"),
("000000","111111","000000","010111","010111","010111","010111","010111","010111","010111","010111","000000","111111","111111","111000","111000","111000","111000","010111","000000","000000","000000","000000","000000","000000","111000","111000","111000","010111","000000","000000","000000","010111","111000","111111","111111","111111","111111","111111","111111","010111","000000","000000","000000","000000","000000","000000","000000","000000","010111","111000","111000","000000","000000","000000","000000"),
("010111","010111","000000","010111","010111","010111","010111","010111","010111","010111","010111","010111","000000","000000","111111","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000","010111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","010111","000000","000000","000000","000000","000000","000000","111000","111000","111000","111000","000000","000000","000000"),
("000000","010111","010111","000000","010111","010111","010111","010111","010111","010111","010111","000000","000000","000000","000000","010111","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","010111","000000","000000","000000","000000","111111","111111","111111","111111","111111","010111","000000","000000","000000","010111","111111","111111","111111","010111","000000","000000","010111","111000","111000","111000","111000","111000","000000","000000","000000"),
("000000","111111","010111","010111","000000","000000","000000","010111","010111","000000","000000","000000","000000","000000","111000","010111","000000","000000","010111","111000","111000","111000","111000","111000","010111","000000","000000","000000","000000","000000","000000","111111","111111","111111","000000","000000","010111","111111","111111","010111","000000","000000","010111","111111","111111","000000","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000"),
("000000","000000","010111","111111","111111","010111","010111","000000","000000","000000","000000","000000","000000","000000","111111","111000","111000","111000","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","111111","111111","000000","010111","010111","010111","010111","010111","000000","010111","010111","000000","010111","111111","111111","000000","111000","111000","111000","111000","111000","111000","000000","000000","000000"),
("000000","000000","000000","111111","000000","010111","010111","000000","000000","000000","000000","000000","000000","000000","010111","111111","111111","111000","111000","111000","010111","010111","000000","000000","000000","000000","000000","000000","000000","000000","111000","111111","000000","010111","000000","111111","111111","111111","010111","010111","010111","000000","010111","000000","111111","111111","000000","111000","111000","111000","111000","111000","111000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","111000","111111","111111","111111","111000","111000","111000","111000","111000","111000","111000","111000","111000","010111","000000","111000","111111","000000","000000","010111","000000","000000","000000","000000","010111","111111","010111","000000","010111","000000","111111","111111","010111","111000","111000","111000","111000","111000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","010111","010111","000000","010111","111111","111111","111111","111111","111000","111111","111000","111000","111000","111000","111000","111000","000000","111000","000000","010111","010111","010111","010111","010111","010111","010111","000000","000000","010111","010111","000000","000000","111111","111111","000000","111000","111000","111000","111000","111000","010111","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","010111","010111","010111","000000","111111","010111","111000","111111","111111","111111","111000","111111","111000","111000","111000","111000","111000","000000","111000","000000","010111","010111","010111","010111","010111","010111","010111","010111","010111","000000","010111","010111","000000","010111","111111","111111","000000","111000","111000","111000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","010111","010111","010111","000000","111111","010111","010111","111111","111000","111111","111000","111000","111000","111000","111000","111000","111000","000000","111111","111111","111111","010111","010111","010111","111111","000000","010111","010111","010111","000000","000000","000000","010111","111111","111111","111111","000000","000000","111000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","010111","010111","010111","000000","111000","111111","111111","010111","010111","010111","111111","111000","111000","111000","111000","010111","010111","000000","111111","111111","111111","010111","010111","111111","111111","111111","000000","010111","010111","000000","000000","000000","000000","000000","010111","111111","111111","111111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","010111","010111","010111","010111","000000","111111","111111","111111","111111","111111","010111","010111","010111","010111","010111","111111","111000","000000","111000","111111","000000","010111","000000","111000","111111","111000","000000","010111","010111","010111","000000","000000","010111","010111","010111","000000","111111","111000","111111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","010111","010111","010111","010111","010111","010111","000000","111000","111111","111111","111111","111111","111111","111111","111000","111000","111000","111000","000000","000000","111000","000000","010111","000000","111000","111000","000000","010111","010111","010111","010111","000000","000000","010111","010111","010111","010111","000000","111111","111000","111000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","010111","010111","010111","010111","010111","010111","000000","000000","111000","111111","111111","111000","111111","111000","111111","111000","111000","111000","111000","000000","000000","000000","010111","010111","000000","000000","010111","000000","111000","010111","000000","000000","010111","010111","010111","010111","010111","000000","000000","111111","111000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","010111","010111","010111","010111","010111","000000","000000","010111","000000","000000","111000","111111","111000","111111","111000","111000","111000","111000","111000","111000","000000","010111","010111","010111","010111","010111","000000","111000","111111","111111","000000","000000","010111","010111","010111","010111","010111","000000","000000","111000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","010111","010111","010111","000000","000000","010111","000000","010111","000000","000000","000000","010111","111000","111111","111000","111000","111000","111000","111000","111000","000000","000000","010111","010111","010111","000000","111000","111000","000000","000000","010111","010111","010111","010111","010111","010111","000000","000000","000000","000000","010111","010111","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","010111","000000","010111","000000","000000","000000","000000","010111","111000","000000","111000","000000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","010111","010111","010111","010111","010111","010111","010111","000000","000000","000000","000000","000000","000000","010111"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","000000","010111","010111","010111","010111","000000","010111","000000","010111","000000","010111","000000","000000","000000","111000","000000","111000","000000","111000","000000","000000","000000","000000","000000","010111","010111","000000","010111","010111","010111","010111","010111","010111","010111","000000","010111","000000","000000","000000","000000","010111","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","111111","111111","111111","000000","000000","010111","000000","010111","000000","010111","000000","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","010111","010111","010111","000000","010111","010111","010111","010111","010111","000000","010111","000000","000000","010111","010111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","111111","111111","111111","111111","111000","111000","000000","000000","111000","111000","000000","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","010111","010111","010111","010111","000000","000000","000000","000000","000000","010111","000000","010111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","111111","111111","111111","111000","111000","111000","000000","000000","111111","111111","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","111000","111000","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","010111","010111","010111","000000","000000","000000","010111","010111","010111","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","111000","111000","000000","000000","010111","000000","111111","111111","111000","000000","010111","000000","000000","111000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","111111","111000","111000","111000","000000","000000","111111","111111","111111","111000","111000","000000","000000","111000","111000","111000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111000","111000","111000","000000","111000","111000","111111","111111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","111111","111111","111111","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"));

Constant HpString : Hp :=( ("000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000110","000110","000110","000110","010110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111000","111000","101001","101001","011010","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","011010","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","111000","101001","101001","011001","010110","010110","010110","000110","000110","000110","000110","000110","000110","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","101011","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","101011","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101011","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000110","000110","000110","000110","010110","101001","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000110","000110","000110","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","011010","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000110","000110","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","011010","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","010110","010110","101010","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000110","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","011010","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","000110","000110","000110","000110","011010","010110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","010110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","101001","111100","111100","111000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","010110","010110","010110","010110","000110","000110","000110","000110","000110","000110","011010","101011","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","010110","000110","000110","000110","000110","011010","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","011010","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","000110","000110","010110","101001","010110","000110","000110","000110","000110","000110","101010","111111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","111100","111100","111100","111100","111100","011001","000110","000110","000110","010110","111111","111111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","101001","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","101010","111111","111111","000000","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","011010","111100","111100","111100","111100","111100","111100","111100","111100","111100","011001","000110","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","000000","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","111100","111100","111100","111100","111000","111100","111100","111100","111100","111000","000110","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","011010","111111","111111","111111","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","011010","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","101001","111100","111100","111000","111000","111100","111100","111100","111100","111100","000110","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","010110","010110","000110","111100","111100","111100","111100","111100","111100","000110","111000","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","000110","010110","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","101011","111111","111111","111111","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","101001","111000","111100","111100","111100","111100","111100","111100","111000","000110","000110","010110","111000","111100","111100","111100","011010","000110","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","011010","111111","111111","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","111100","101000","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","000110","000110","000110","010110","101001","011010","010110","000110","000110","000110","000110","101010","111111","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","000110","000110","000110","101001","111100","111100","111100","111100","101001","000110","000110","000110","000110","101011","111111","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","011010","111111","111111","000000"),
("000000","000000","000000","000110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","010110","111111","111111","111111"),
("000000","000000","000000","000110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","010110","111111","111111","111111"),
("000000","000000","000000","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","011010","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","010110","111111","111111","111111"),
("000000","000000","000000","000000","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","011010","101011","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","011010","111111","111111","111111"),
("000000","000000","000000","000000","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","011010","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","010110","101011","111111","011010","000110","000110","000110","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","101010","111111","111111","111111"),
("000000","000000","000000","000000","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","011001","000110","000110","000110","000110","000110","010110","101011","111111","111111","101010","000110","000110","000110","000110","101001","111100","111100","111100","101001","000110","000110","000110","010110","111111","111111","111111","111111"),
("000000","000000","000000","000000","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","000110","000110","000110","000110","011010","101011","111111","111111","111111","111111","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","101010","111111","111111","111111","111111"),
("000000","000000","000000","000000","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","000110","010110","101010","111111","111111","111111","111111","111111","111111","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","101010","111111","111111","111111","111111","000000"),
("000000","000000","000000","000000","000110","000110","000110","011010","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","011010","101010","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000110","010110","000110","000110","000110","000110","000110","010110","101010","111111","111111","111111","111111","111111","000000"),
("000000","000000","000000","000000","000110","000110","000110","010110","101001","101001","101001","101001","101001","101001","101001","101001","010110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","011010","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","111111","101011","101010","101010","101010","101011","111111","111111","111111","111111","111111","111111","000000","000000"),
("000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","011010","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","011010","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","011010","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000110","000110","010110","010110","010110","010110","010110","010110","010110","010110","010110","010110","011010","000110","000110","000110","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","010110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","101010","000110","000110","000110","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","010110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","101010","000110","000110","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","011010","101010","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","101010","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","011010","101001","101001","101001","101001","101001","101001","101001","011010","000110","000110","000110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","010110","010110","010110","010110","010110","010110","010110","010110","010110","011010","101011","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000")); 

Constant AtString : At :=( ("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","101011","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","101010","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","010110","101001","000110","000110","000110","101010","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","101010","111111","111111","000000","000110","000110","000110","000110","000110","000110","000110","010110","111000","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","010110","000110","000110","010110","111111","111111","011010","000110","000110","000110","000110","000110","010110","111000","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","101001","111100","101001","000110","000110","000110","101010","111111","011010","000110","000110","000110","011010","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","000110","000110","000110","011010","111111","011010","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","101001","111100","111100","111100","101001","000110","000110","000110","101011","011010","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","000110","000110","000110","101010","101010","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","010110","000110","000110","000110","101010","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","011010","011010","011010","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","000110","000110","000110","000110","000110","101010","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","010110","010110","010110","010110","000110","000110","000110","101010","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","011010","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","011010","111111","111111","111111","000000","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","011010","111111","111111","111111","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","011010","111111","111111","011010","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","011010","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","011010","111111","101010","000110","000110","000110","000110","010110","101001","010110","000110","000110","000110","000110","000110","101010","111111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","011010","101010","011010","000110","000110","000110","111100","111100","111100","111100","111100","011001","000110","000110","000110","010110","111111","111111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","101001","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","101010","111111","111111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","101000","101001","111100","111100","111100","111100","111100","111100","111100","101001","011001","011001","111100","111100","111100","111100","111100","111100","111100","111000","011001","011001","011001","011001","011001","000110","000110","000110","000110","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","011010","111111","111111","111111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","011001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","000110","000110","000110","010110","111000","101001","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","011010","000110","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","000110","000110","101001","111100","111100","111100","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","011010","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","010110","111100","111100","111100","111100","111100","010110","000110","000110","010110","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","101011","111111","111111","111111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","010110","111000","111100","111100","111100","011010","000110","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000110","000110","000110","000110","011010","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","101001","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","011010","111111","111111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","111100","111000","111100","111100","111100","111100","111100","111100","111100","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","000110","000110","000110","000110","010110","101001","011010","010110","000110","000110","000110","000110","101010","111111","000000","000000","000000"),
("000000","000000","000000","000000","000110","000110","000110","000110","011010","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","101000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","000110","000110","000110","101001","111100","111100","111100","111100","101001","000110","000110","000110","000110","101011","111111","000000","000000"),
("000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","011010","111111","111111","000000"),
("000000","000000","000000","000110","000110","000110","000110","011010","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","010110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","010110","111111","111111","111111"),
("000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","101010","011010","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","010110","111111","111111","111111"),
("000000","000000","000110","000110","000110","000110","011010","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","101011","101010","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","010110","111111","111111","111111"),
("000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","101010","111111","111111","010110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","011001","101000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","010110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","011010","111111","111111","111111"),
("000000","000110","000110","000110","000110","011010","111100","111100","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","000110","101011","111111","111111","101010","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","111100","000110","011001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","011001","000110","000110","000110","000110","101010","011010","000110","000110","000110","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","101010","111111","111111","111111"),
("000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","011010","111111","111111","111111","101011","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","101001","111000","111100","111100","111100","111100","101001","010110","000110","000110","000110","000110","000110","101010","111111","101010","000110","000110","000110","000110","101001","111100","111100","111100","101001","000110","000110","000110","010110","111111","111111","111111","111111"),
("000110","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","011001","000110","000110","000110","101011","111111","111111","111111","111111","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","101010","111111","111111","111111","011010","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","101010","111111","111111","111111","111111"),
("000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","011010","111111","111111","111111","111111","000000","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","011010","101010","111111","111111","111111","111111","111111","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","101010","111111","111111","111111","111111","000000"),
("000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","101010","111111","111111","111111","111111","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","011001","000110","000110","000110","000110","000110","000110","000110","000110","010110","011010","101011","111111","111111","111111","111111","111111","111111","000000","000000","000110","010110","000110","000110","000110","000110","000110","010110","101010","111111","111111","111111","111111","111111","000000"),
("000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","011010","111111","111111","111111","111111","000000","000000","000000","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","011010","101010","101010","101010","101011","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","111111","101011","101010","101010","101010","101011","111111","111111","111111","111111","111111","111111","000000","000000"),
("000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","101010","111111","111111","111111","111111","000000","000000","000000","000000","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","010110","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000"),
("000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","111111","111111","111111","111111","000000","000000","000000","000000","000000","000110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","101010","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000"),
("000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","011010","101011","111111","111111","111111","111111","000000","000000","000000","000000","000000","000110","000110","000110","000110","011010","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000110","101010","101010","101010","101010","101010","101010","101010","101010","101010","101010","101010","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111000","101001","101001","011001","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","101011","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","101010","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","011010","101010","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","101010","101010","101010","101010","101011","101011","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"));

Constant DefString : Def :=( ("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010110","000110","000110","000110","000110","000110","000110","000110","101010","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","000110","000110","000110","000110","000110","000110","011010","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","101001","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","000110","101010","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","011010","111000","111100","111100","111100","111100","111100","111100","111100","111000","010110","000110","000110","000110","000110","101010","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000110","000110","000110","000110","000110","000110","010110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","000110","011010","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","000110","101011","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","000110","101010","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","011010","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","101010","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","010110","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","011010","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","010110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","101010","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000110","000110","000110","011010","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","011010","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","000110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","010110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","101001","111000","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","101010","111111","111111","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","010110","111100","111100","111100","111100","101001","000110","000110","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","101011","101010","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","011001","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","011010","111100","111000","010110","000110","000110","000110","000110","000110","101010","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","011010","000110","000110","000110","000110","000110","011010","101011","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","111100","111000","101001","101001","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","000110","000110","000110","000110","000110","010110","101010","101011","101010","011010","010110","010110","011010","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000110","000110","000110","000110","111100","101001","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","011001","000110","000110","010110","101011","101010","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000110","000110","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","011001","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","010110","101010","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","011010","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","011010","111100","111100","111100","111100","111100","111100","111100","111000","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","010110","000110","000110","000110","000110","010110","101001","010110","000110","000110","000110","000110","000110","101010","111111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","011001","111100","111100","111100","111100","111100","111100","111100","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","000110","000110","111100","111100","111100","111100","111100","011001","000110","000110","000110","010110","111111","111111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","101010","111111","111111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","011010","111111","111111","111111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","011010","000110","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","101001","111100","111100","111100","111100","111100","111100","011010","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","101001","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","011010","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","101011","111111","111111","111111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","101001","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","111100","111100","111100","111100","111100","111100","101000","101001","111100","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","000110","000110","000110","101010","011010","000110","000110","000110","010110","111000","111100","111100","111100","011010","000110","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","111100","111100","111000","000110","111000","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","101010","101010","101011","111111","101011","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","011010","111111","111111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","111100","111100","111100","111100","101001","111000","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","101011","111111","111111","111111","111111","101011","010110","000110","000110","000110","000110","000110","010110","101001","011010","010110","000110","000110","000110","000110","101010","111111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","111100","111100","111100","111100","111100","111100","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101011","111111","111111","111111","111111","111111","000110","000110","000110","000110","000110","101001","111100","111100","111100","111100","101001","000110","000110","000110","000110","101011","111111","000000","000000"),
("000000","000000","000000","000000","000000","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","011010","111111","111111","000000"),
("000000","000000","000000","000000","000000","000000","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","011001","011010","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","010110","111111","111111","111111"),
("000000","000000","000000","000000","000000","000000","000110","000110","000110","011010","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","011001","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","010110","111111","111111","111111"),
("000000","000000","000000","000000","000000","000000","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","010110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","010110","111111","111111","111111"),
("000000","000000","000000","000000","000000","000000","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","011010","000110","000110","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","010110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","011010","111111","111111","111111"),
("000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111000","101001","011010","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","011010","000110","000110","011010","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","101010","111111","111111","111111"),
("000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","011001","010110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","011010","011010","000110","000110","000110","000110","010110","101001","111000","111100","111100","111100","111100","111000","101001","011010","010110","000110","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000","000110","000110","000110","000110","000110","101001","111100","111100","111100","101001","000110","000110","000110","010110","111111","111111","111111","111111"),
("000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","011010","101011","111111","111111","011010","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","101010","111111","111111","111111","111111"),
("000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","011010","101010","101010","101111","111111","111111","111111","111111","111111","101010","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","101010","111111","111111","111111","111111","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","010110","011010","101010","101010","101011","101011","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000110","101010","010110","000110","000110","000110","000110","000110","000110","000110","000110","010110","011010","101010","011010","000110","000110","010110","111100","111100","111100","111100","111100","111100","111000","111000","101001","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000","000000","000000","000000","000110","010110","000110","000110","000110","000110","000110","010110","101010","111111","111111","111111","111111","111111","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","111111","101011","101010","101010","101010","101010","101010","101010","101011","111111","111111","111111","101010","000110","000110","000110","101001","011010","010110","010110","000110","000110","000110","000110","000110","000110","000110","000110","101011","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","111111","101011","101010","101010","101010","101011","111111","111111","111111","111111","111111","111111","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","101011","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","101010","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","101010","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","010110","010110","011010","101010","101010","101010","101011","101011","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"));

Constant SpString : Sp :=( ("000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","010110","010110","010110","010110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000110","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","011010","000110","000110","000110","000110","000110","000110","010110","101011","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000110","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","011010","000110","000110","000110","000110","101010","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000110","000110","000110","011001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","011001","000110","000110","000110","101010","101011","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","000110","000110","010110","101011","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111000","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","000110","000110","000110","011010","010110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000110","000110","000110","011010","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","000110","010110","101001","111000","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","010110","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","000110","000110","010110","101001","111100","111100","111100","111100","111100","000110","101001","111100","111100","111000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111000","000110","010110","010110","010110","010110","000110","000110","000110","000110","000110","000110","011010","101011","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000110","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","000110","000110","000110","011010","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","010110","000110","000110","000110","000110","011010","000110","000110","000110","000110","000110","000110","000110","000110","000110","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","011010","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","000110","000110","010110","101001","010110","000110","000110","000110","000110","000110","101010","111111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000110","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","111100","111100","111100","111100","111100","011001","000110","000110","000110","010110","111111","111111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000110","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","101001","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","101010","111111","111111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","011010","111100","111100","111100","111100","111100","111100","111100","111100","111100","011001","000110","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","000000","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","111100","111100","111100","111100","111000","111100","111100","111100","111100","111000","000110","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","011010","111111","111111","111111","000000","000000","000000"),
("000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","101001","111100","111100","111000","111000","111100","111100","111100","111100","111100","000110","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000"),
("000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","010110","010110","000110","111100","111100","111100","111100","111100","111100","000110","111000","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000"),
("000000","000000","000110","000110","000110","000110","111100","111100","010110","000110","000110","000110","000110","000110","000110","000110","011001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","000110","010110","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","101011","111111","111111","111111","000000","000000","000000"),
("000000","000000","000110","000110","000110","010110","111100","111100","111100","111000","010110","000110","000110","000110","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","101001","111000","111100","111100","111100","111100","111100","111100","111000","000110","000110","010110","111000","111100","111100","111100","011010","000110","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000"),
("000000","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","101001","010110","000110","000110","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","011010","111111","111111","000000","000000","000000"),
("000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","011001","010110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","000110","000110","000110","010110","101001","011010","010110","000110","000110","000110","000110","101010","111111","000000","000000","000000"),
("000000","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","000110","000110","000110","101001","111100","111100","111100","111100","101001","000110","000110","000110","000110","101011","111111","000000","000000"),
("000110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","011010","111111","111111","000000"),
("000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","000110","000110","000110","111000","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","010110","111111","111111","111111"),
("000110","000110","000110","011010","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","010110","111111","111111","111111"),
("000110","000110","000110","010110","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","011010","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","010110","111111","111111","111111"),
("000110","000110","000110","000110","000110","000110","011010","111000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","011010","101011","000110","000110","000110","101001","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","011010","111111","111111","111111"),
("000110","000110","000110","000110","000110","000110","000110","000110","000110","011010","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","000110","010110","101011","111111","011010","000110","000110","000110","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","101010","111111","111111","111111"),
("000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","011010","101001","111000","111100","111100","111100","111100","111100","101001","010110","000110","101001","111100","111100","111100","111100","111100","111100","111100","111100","111100","111000","011001","000110","000110","000110","000110","000110","010110","101011","111111","111111","101010","000110","000110","000110","000110","101001","111100","111100","111100","101001","000110","000110","000110","010110","111111","111111","111111","111111"),
("000000","000000","000000","101010","101010","011010","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","011001","111100","111100","111100","111100","111100","111100","111100","111100","000110","000110","000110","000110","000110","000110","000110","011010","101011","111111","111111","111111","111111","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","101010","111111","111111","111111","111111"),
("000000","000000","000000","000000","111111","111111","101111","101010","011010","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","011010","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","000110","000110","010110","101010","111111","111111","111111","111111","111111","111111","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","101010","111111","111111","111111","111111","000000"),
("000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","101011","101010","011010","010110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","011010","101010","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000110","010110","000110","000110","000110","000110","000110","010110","101010","111111","111111","111111","111111","111111","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","101011","101011","101010","101010","101010","101010","101010","011010","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","011010","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","111111","101011","101010","101010","101010","101011","111111","111111","111111","111111","111111","111111","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","011010","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","010110","000110","000110","011010","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","011010","000110","000110","010110","111100","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","011010","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","011010","000110","000110","010110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","010110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","101001","000110","000110","000110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","111100","111100","111100","111100","111100","111100","111100","111100","111000","000110","000110","000110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","011010","101001","101001","101001","101001","101001","101001","101001","011010","000110","000110","000110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","010110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","000110","101010","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000110","000110","010110","010110","010110","010110","010110","010110","010110","010110","010110","011010","101011","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"));


constant FireblastString : Fireblast :=(('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','1','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','1','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','0','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','1','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','1','1','1','1','1','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','1','1','1','1','1','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','0','0','1','1','1','1','0','0','0','0','0','1','1','1','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','1','0','1','1','1','1','0','0','0','0','0','1','1','1','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','1','1','1','1','0','0','0','0','0','1','1','1','0','0','1','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','1','1','1','1','0','0','0','0','0','1','1','1','1','0','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','1','1','1','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','1','1','1','0','0','1','1','1','1','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','0','0','1','1','1','1','1','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','1','1','1','0','0','0','1','1','1','1','1','0','0','1','1','0','0','0','1','1','1','1','0','0','0','1','1','1','1','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));





constant LeafBladeString : LeafBlade :=(('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','0','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','1','1','1','0','0','0','0','0','1','1','1','1','0','0','1','1','1','0','0','0','0','0','1','1','1','1','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','0','1','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','1','1','1','0','0','0','0','0','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','0','0','0','0','0','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','1','1','1','1','0','0','1','1','1','0','0','0','0','0','1','1','1','1','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','1','1','1','1','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','0','0','0','0','0','1','1','1','1','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','0','0','1','1','1','0','0','0','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','0','1','1','1','1','0','0','1','1','1','0','0','0','1','1','1','1','1','0','0','1','1','1','1','0','0','0','1','1','1','1','1','0','0','0','1','1','1','1','0','0','0','0','1','1','0','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','1','0','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','0','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));



constant MegaPunchString : Megapunch:=(('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','1','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','1','1','1','0','1','1','1','0','0','0','0','0','1','1','1','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','1','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','0','1','1','1','1','1','0','0','0','1','1','1','0','0','0'),
('0','0','0','1','1','1','0','1','1','1','1','0','0','0','0','1','1','1','0','1','1','1','0','0','0','1','1','1','1','0','0','0','0','1','1','1','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0'),
('0','0','0','1','1','1','0','0','1','1','1','0','0','0','1','1','1','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','1','1','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0'),
('0','0','0','1','1','1','0','0','1','1','1','0','0','0','1','1','1','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','1','1','1','0','0','0','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0'),
('0','0','0','1','1','1','0','0','1','1','1','1','0','1','1','1','1','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0'),
('0','0','0','1','1','1','0','0','0','1','1','1','0','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0'),
('0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0'),
('0','0','0','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0'),
('0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','0','0','1','1','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','1','1','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','1','1','1','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0'),
('0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));


constant SurfString: Surf:=(('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0'),
('0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0','0'),
('0','0','0','0','1','1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','0'),
('0','0','0','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0'),
('0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
('0','0','0','1','1','1','1','1','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0'),
('0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','1','1','1','1','1','1','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','1','1','1','1','1','0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','1','1','1','0','0','0','0','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0'),
('0','0','1','1','1','1','0','0','0','1','1','1','1','0','0','0','1','1','1','1','0','0','1','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0'),
('0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','1','1','1','0','0','1','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0'),
('0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','1','0','1','1','1','0','0','1','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));



constant AustossBackString : Pokemon :=(("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","010001","111111","111111","100111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","111111","111111","111111","100111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","100111","111111","111111","100111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","000000","111111","111111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","010001","100111","100111","111111","111111","100111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100111","111111","111111","111111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","100111","100111","111111","111111","100111","100111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","100111","111111","111111","100111","100111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","100111","100111","111111","111111","100111","100111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","100111","111111","111111","100111","100111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","010001","100111","100111","100111","111111","111111","100111","100111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","000000","111111","111111","100111","000000","000000","000000","000000","000000","010001","000000","000000","000000","000000","100111","111111","111111","100111","100111","100111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100111","100111","100111","111111","111111","111111","100111","100111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","100111","100111","100111","000000","000000","000000","000000","111111","111111","100111","000000","100111","111111","100111","100111","100111","010001","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100111","100111","100111","111111","000000","000000","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","100111","100111","010001","000000","000000","000000","000000","000000","111111","111111","100111","000000","100111","100111","100111","100111","100111","010001","010001","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","100111","100111","100111","000000","010001","010001","000000","010001","000000","000000","000000","000000","000000","000000","000000","000000","111111","100111","100111","010001","000000","000000","000000","000000","000000","100111","100111","100111","100111","000000","100111","111111","100111","100111","100111","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","100111","000000","010001","010001","100111","100111","100111","000000","000000","000000","000000","000000","000000","100111","100111","100111","000000","000000","000000","000000","000000","000000","100111","100111","100111","010001","000000","111111","111111","100111","100111","010001","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","010001","010001","100111","010001","100111","010001","100111","000000","000000","000000","000000","100111","100111","100111","010001","000000","000000","000000","010001","100111","100111","100111","100111","010001","111111","111111","111111","100111","010001","010001","010001","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","100111","010001","100111","010001","010001","000000","000000","100111","100111","100111","000000","000000","000000","000000","100111","111111","111111","100111","100111","100111","000000","111111","111111","010001","010001","010001","010001","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","100111","010001","000000","000000","100111","100111","100111","010001","000000","000000","000000","100111","111111","111111","111111","100111","100111","100111","000000","100111","100111","010001","010001","010001","010001","010001","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","000000","000000","100111","100111","100111","100111","000000","000000","000000","100111","111111","111111","100111","100111","100111","100111","100111","000000","000000","100111","100111","010001","010001","010001","010001","010001","010001","000000","100111","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","100111","100111","100111","100111","010001","000000","000000","000000","111111","111111","111111","100111","111111","100111","100111","010001","000000","111111","111111","000000","010001","010001","100111","010001","100111","010001","000000","100111","100111","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100111","100111","100111","010001","000000","000000","000000","111111","111111","111111","100111","111111","100111","100111","100111","100111","111111","111111","100111","010001","000000","010001","010001","100111","010001","000000","100111","000000","100111","100111","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","100111","100111","100111","000000","000000","000000","100111","111111","111111","111111","100111","111111","100111","100111","100111","100111","100111","100111","100111","010001","010001","010001","000000","100111","010001","000000","100111","100111","000000","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","100111","010001","000000","000000","100111","111111","100111","111111","100111","100111","100111","100111","100111","100111","100111","100111","100111","010001","010001","010001","000000","010001","000000","000000","100111","100111","100111","000000","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010001","010001","010001","000000","000000","100111","111111","100111","111111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","010001","010001","010001","000000","010001","010001","010001","100111","100111","000000","100111","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","010001","000000","000000","000000","000000","000000","010001","010001","010001","010001","000000","000000","100111","111111","100111","111111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","010001","100111","010001","010001","010001","010001","010001","100111","010001","100111","010001","100111","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","010001","111111","111111","000000","000000","010001","000000","000000","000000","000000","010001","000000","100111","111111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","010001","100111","010001","010001","010001","010001","010001","010001","010001","100111","100111","100111","100111","100111","100111","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","000000","111111","111111","000000","100111","010001","000000","000000","000000","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","010001","100111","010001","100111","010001","010001","010001","100111","010001","100111","100111","100111","100111","100111","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","010001","111111","100111","000000","000000","000000","111111","111111","000000","010001","100111","010001","100111","010001","000000","100111","100111","100111","100111","010001","000000","100111","100111","100111","010001","000000","000000","000000","100111","010001","100111","010001","100111","010001","100111","010001","100111","100111","100111","100111","100111","100111","100111","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","100111","111111","000000","000000","000000","010001","100111","111111","000000","010001","100111","010001","100111","000000","100111","100111","010001","000000","111111","100111","000000","000000","000000","100111","100111","100111","100111","000000","100111","010001","100111","010001","100111","010001","100111","010001","100111","100111","100111","100111","100111","100111","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","010001","000000","000000","000000","000000","111111","100111","000000","100111","010001","100111","010001","010001","000000","000000","100111","111111","111111","111111","111111","111111","100111","100111","100111","100111","100111","100111","100111","100111","010001","100111","010001","100111","010001","100111","100111","100111","100111","100111","100111","100111","100111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","010001","100111","100111","000000","000000","000000","000000","000000","010001","111111","100111","000000","010001","010001","010001","010001","000000","100111","100111","111111","111111","111111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","000000","010001","100111","100111","100111","100111","100111","100111","100111","100111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","100111","010001","000000","000000","000000","000000","000000","000000","100111","100111","000000","010001","010001","010001","010001","010001","000000","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","111111","111111","100111","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","010001","100111","100111","000000","000000","000000","000000","000000","000000","000000","100111","100111","000000","010001","010001","010001","010001","010001","000000","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","100111","111111","111111","111111","111111","100111","111111","100111","111111","100111","100111","010001","010001","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","100111","100111","000000","000000","000000","000000","000000","000000","000000","100111","100111","010001","010001","010001","010001","010001","010001","000000","100111","010001","100111","100111","100111","100111","100111","100111","100111","010001","100111","100111","100111","100111","100111","111111","111111","111111","100111","111111","100111","111111","100111","100111","000000","010001","010001","010001","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","100111","100111","000000","000000","000000","000000","000000","010001","100111","000000","010001","010001","000000","010001","000000","010001","000000","010001","100111","010001","100111","010001","100111","010001","100111","010001","100111","010001","100111","100111","100111","100111","100111","111111","100111","111111","100111","100111","100111","100111","100111","010001","010001","010001","010001","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","100111","010001","000000","000000","000000","000000","100111","100111","010001","010001","000000","010001","000000","010001","000000","010001","010001","010001","100111","010001","100111","010001","100111","010001","000000","010001","100111","010001","100111","100111","100111","100111","100111","100111","100111","100111","100111","010001","010001","010001","000000","010001","010001","010001","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","100111","100111","000000","000000","000000","010001","100111","000000","010001","010001","010001","000000","010001","000000","010001","010001","010001","010001","010001","100111","010001","100111","000000","010001","010001","100111","010001","100111","010001","100111","100111","100111","100111","010001","010001","010001","010001","010001","010001","010001","010001","010001","010001","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","100111","010001","000000","000000","000000","100111","100111","010001","010001","010001","010001","010001","010001","000000","010001","010001","010001","010001","010001","010001","010001","010001","100111","010001","100111","010001","100111","010001","100111","010001","010001","010001","010001","010001","010001","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","100111","000000","000000","000000","010001","100111","000000","010001","010001","010001","010001","010001","010001","010001","000000","010001","010001","010001","010001","100111","010001","100111","010001","100111","010001","100111","010001","010001","010001","010001","010001","010001","010001","010001","000000","000000","000000","100111","010001","100111","010001","100111","010001","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","010001","100111","100111","000000","000000","000000","100111","100111","000000","010001","010001","010001","010001","010001","010001","010001","000000","010001","010001","010001","010001","010001","100111","010001","100111","010001","100111","010001","100111","010001","010001","010001","010001","010001","010001","000000","100111","010001","100111","010001","100111","010001","100111","010001","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","100111","100111","000000","000000","000000","100111","100111","000000","010001","010001","010001","010001","100111","010001","100111","010001","010001","010001","010001","010001","010001","000000","000000","010001","100111","010001","100111","010001","010001","010001","010001","010001","010001","000000","100111","010001","100111","010001","100111","010001","010001","010001","010001","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","100111","100111","000000","000000","000000","010001","100111","100111","010001","100111","010001","100111","010001","100111","010001","010001","000000","010001","010001","010001","000000","100111","100111","000000","000000","100111","010001","100111","010001","010001","010001","010001","010001","010001","010001","100111","010001","010001","010001","010001","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","100111","100111","000000","000000","000000","000000","100111","100111","000000","010001","100111","010001","100111","010001","100111","010001","000000","010001","000000","000000","100111","100111","100111","100111","100111","000000","000000","000000","010001","010001","010001","010001","010001","010001","010001","010001","010001","010001","010001","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","100111","100111","010001","000000","000000","000000","000000","100111","100111","000000","100111","010001","100111","010001","100111","010001","010001","000000","010001","100111","010001","100111","010001","100111","010001","100111","100111","010001","010001","010001","010001","010001","010001","010001","010001","010001","010001","010001","010001","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","100111","100111","000000","000000","000000","000000","000000","010001","100111","100111","010001","100111","010001","100111","010001","010001","010001","010001","000000","010001","100111","010001","100111","010001","100111","010001","010001","010001","010001","010001","010001","010001","010001","010001","010001","010001","000000","010001","000000","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","100111","100111","000000","000000","000000","000000","000000","000000","100111","100111","000000","010001","010001","010001","010001","010001","000000","010001","000000","010001","010001","100111","010001","100111","010001","010001","010001","010001","010001","010001","010001","000000","010001","000000","010001","000000","010001","000000","010001","000000","010001","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","100111","100111","000000","000000","000000","000000","000000","000000","100111","100111","000000","010001","010001","010001","010001","000000","010001","000000","000000","010001","010001","010001","010001","010001","010001","010001","010001","010001","010001","000000","000000","010001","000000","010001","000000","010001","000000","010001","000000","010001","000000","010001","000000","000000","000000","000000","000000","000000","000000","000000","000000"));

constant BisaflorBackString : Pokemon :=(("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110110","000000","000000","111111","111111","110110","110110","110110","000000","000000","000000","000000","000000","000000","110110","000000","111111","111111","111111","110110","110110","110110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110110","000000","000000","111111","110110","110110","110110","111111","111111","111111","110110","110110","110110","110110","000000","000000","110110","111111","111111","111111","110110","110110","110110","111111","111111","111111","110110","110110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","110110","111111","110110","111111","110110","110110","110110","111111","111111","111111","110110","110110","110110","110110","000000","000000","111111","110110","110110","110110","110110","111111","111111","111111","110110","110110","110110","110110","110110","110110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110110","111111","110110","111111","110110","111111","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","000000","000000","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","000000","110110","000000","000000","110110","110110","110110","110110","110110","110110","110110","110110","110110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","110110","000000","111111","110110","111111","110110","111111","110110","111111","000000","000000","000000","000000","110110","110110","110110","110110","110110","000000","000000","111111","000000","000000","111111","000000","000000","110110","110110","110110","110110","000000","000000","000000","110110","110110","110110","110110","110110","110110","110110","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","111111","110110","111111","111111","111111","111111","111111","110110","110110","111111","111111","110110","000000","000000","110110","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","110110","000000","110110","110110","110110","110110","110110","110110","110110","111111","111111","111111","110110","110110","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","110110","111111","110110","110110","111111","111111","111111","111111","111111","110110","110110","110110","110110","110110","110110","110110","110110","000000","111111","000000","111111","110110","000000","000000","000000","000000","110110","111111","000000","111111","000000","110110","110110","110110","110110","110110","110110","110110","111111","111111","111111","110110","110110","110110","110110","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","110110","110110","111111","110110","111111","110110","111111","110110","111111","110110","110110","110110","110110","110110","110110","110110","000000","111111","111111","000000","000000","111111","111111","111111","111111","000000","000000","111111","111111","000000","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","110110","111111","110110","111111","110110","111111","110110","111111","110110","110110","110110","110110","110110","110110","110110","110110","000000","111111","111111","000000","111111","000000","111111","111111","000000","111111","000000","111111","000000","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","110110","110110","110110","111111","000000","000000","110110","111111","110110","110110","110110","111111","111111","111111","110110","110110","110110","110110","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","110110","110110","110110","110110","110110","110110","111111","111111","111111","110110","110110","110110","110110","110110","110110","110110","110110","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","110110","110110","000000","000000","111111","110110","111111","110110","111111","110110","111111","111111","111111","110110","110110","110110","110110","110110","000000","000000","111111","000000","000000","000000","000000","000000","111111","000000","110110","110110","110110","110110","110110","110110","111111","111111","111111","111111","111111","110110","110110","110110","110110","110110","110110","110110","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","110110","000000","110110","110110","110110","111111","110110","111111","110110","110110","110110","110110","110110","110110","110110","110110","000000","000000","000000","110110","110110","110110","110110","110110","110110","110110","110110","000000","000000","110110","110110","110110","110110","110110","110110","111111","111111","110110","110110","110110","110110","110110","110110","000000","110110","110110","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","000000","000000","110110","110110","110110","110110","111111","111111","110110","110110","110110","110110","110110","110110","110110","000000","000000","000000","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","000000","110110","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","000000","000000","000000","111111","110110","110110","110110","110110","111111","111111","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","000000","000000","000000","000000","110110","110110","110110","110110","110110","110110","110110","110110","110110","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","110110","110110","110110","110110","110110","110110","110110","110110","000000","000000","000000","000000","111111","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","111111","111111","111111","110110","110110","110110","110110","110110","000000","000000","000000","000000","000000","110110","110110","110110","110110","110110","110110","110110","110110","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","110110","110110","110110","110110","110110","110110","110110","000000","000000","000000","000000","111111","110110","111111","110110","110110","110110","110110","110110","110110","110110","110110","111111","111111","111111","111111","111111","110110","110110","110110","110110","110110","000000","111111","111111","111111","000000","110110","110110","110110","110110","110110","110110","110110","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","110110","110110","110110","110110","110110","000000","000000","000000","000000","111111","110110","111111","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","111111","111111","111111","111111","111111","110110","110110","110110","110110","000000","000000","111111","111111","111111","000000","110110","110110","110110","110110","110110","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","110110","110110","110110","000000","000000","000000","000000","000000","110110","111111","110110","110110","110110","111111","111111","111111","110110","110110","110110","110110","110110","110110","111111","111111","111111","110110","110110","110110","110110","110110","110110","000000","000000","000000","111111","111111","000000","110110","110110","110110","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110110","110110","110110","110110","110110","111111","111111","111111","111111","111111","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","000000","011110","011110","000000","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110110","110110","110110","110110","110110","110110","111111","111111","111111","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","000000","011110","011110","011110","011110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","000000","000000","000000","011110","011110","011110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","000000","011110","011110","000000","000000","011110","011110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","011110","111111","011110","000000","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","000000","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","000000","000000","000000","011110","011110","011110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","011110","111111","011110","111111","011110","000000","110110","110110","110110","110110","110110","110110","110110","110110","110110","000000","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","000000","011110","011110","011110","000000","000000","011110","011110","011110","011110","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","011110","111111","011110","000000","011110","011110","011110","000000","000000","000000","110110","110110","110110","110110","110110","000000","000000","110110","110110","110110","110110","110110","110110","110110","110110","000000","000000","000000","011110","011110","011110","111111","111111","000000","000000","011110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","000000","011110","111111","011110","111111","000000","011110","011110","011110","011110","000000","000000","000000","110110","110110","110110","110110","000000","000000","000000","110110","110110","110110","110110","110110","000000","000000","000000","000000","011110","011110","011110","011110","011110","011110","111111","111111","000000","011110","011110","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","011110","111111","011110","111111","000000","011110","011110","000000","011110","000000","000000","011110","011110","000000","000000","000000","000000","000000","011110","011110","000000","000000","000000","000000","000000","011110","000000","011110","011110","011110","011110","000000","011110","011110","011110","011110","011110","111111","000000","011110","011110","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","011110","000000","011110","011110","011110","000000","011110","011110","000000","000000","011110","111111","011110","011110","011110","011110","111111","000000","011110","011110","011110","011110","000000","000000","000000","011110","011110","011110","000000","011110","011110","011110","000000","011110","011110","011110","011110","011110","011110","011110","111111","011110","011110","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","111111","111111","000000","011110","011110","000000","011110","011110","000000","111111","011110","111111","011110","111111","011110","011110","011110","111111","000000","011110","011110","011110","011110","011110","011110","000000","000000","011110","011110","000000","000000","011110","000000","011110","011110","011110","000000","011110","011110","011110","011110","011110","011110","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","111111","000000","000000","011110","011110","000000","000000","011110","000000","011110","111111","000000","000000","000000","011110","011110","111111","000000","011110","011110","011110","011110","011110","011110","011110","011110","011110","000000","000000","000000","000000","011110","000000","011110","011110","011110","000000","011110","011110","000000","011110","011110","011110","011110","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","111111","011110","000000","011110","011110","011110","000000","000000","000000","011110","000000","000000","111111","011110","111111","011110","011110","111111","000000","011110","011110","011110","011110","000000","000000","011110","011110","011110","011110","000000","000000","000000","000000","000000","011110","011110","000000","011110","011110","011110","000000","011110","011110","011110","011110","011110","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","011110","111111","000000","011110","000000","000000","000000","000000","000000","000000","111111","111111","011110","111111","011110","111111","011110","011110","000000","011110","011110","011110","011110","011110","000000","000000","000000","011110","011110","000000","000000","011110","000000","011110","011110","011110","000000","011110","011110","011110","000000","011110","011110","000000","011110","011110","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","011110","011110","000000","000000","000000","000000","011110","000000","000000","111111","111111","011110","111111","011110","111111","011110","111111","000000","011110","011110","011110","011110","011110","011110","011110","011110","000000","000000","000000","000000","011110","000000","011110","000000","011110","011110","000000","011110","011110","011110","000000","011110","011110","000000","011110","011110","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","011110","000000","000000","111111","000000","011110","000000","011110","000000","011110","011110","111111","000000","000000","011110","011110","111111","000000","011110","011110","011110","000000","000000","011110","011110","011110","011110","011110","000000","011110","000000","011110","000000","011110","000000","000000","000000","011110","011110","000000","011110","011110","011110","000000","011110","011110","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","000000","011110","000000","011110","000000","000000","000000","000000","011110","011110","011110","111111","000000","011110","011110","011110","011110","000000","000000","000000","011110","011110","011110","000000","000000","011110","011110","011110","011110","011110","000000","000000","011110","011110","000000","011110","011110","000000","000000","011110","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","011110","011110","011110","000000","000000","000000","011110","011110","011110","011110","011110","011110","000000","011110","011110","011110","011110","011110","011110","000000","000000","011110","000000","000000","011110","011110","011110","011110","011110","011110","011110","000000","000000","000000","000000","011110","011110","000000","000000","011110","000000","000000","000000","000000","000000","000000"));

constant GallopaBackString : Pokemon :=(("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","111100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111100","111100","111100","111100","111100","111100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111100","110100","111100","111100","111100","111100","111100","110100","000000","000000","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","000000","110100","111100","111100","111100","111100","111100","110100","110100","111100","111100","111100","110100","000000","000000","000000","000000","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111100","111100","111100","111100","111100","110100","110100","111100","111100","111100","110100","000000","000000","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111100","110100","111100","110100","111100","110100","111100","111100","111100","110100","110100","111100","111100","110100","000000","000000","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","000000","000000","000000","000000","000000","000000","110100","110100","111100","110100","111100","110100","111100","111100","111100","110100","111100","110100","111100","110100","110100","110100","000000","000000","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","110100","111100","111100","111100","111100","110100","000000","000000","000000","000000","000000","110100","110100","111100","110100","110100","110100","111100","110100","111100","111100","111100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111100","111100","111100","111100","111100","111100","111100","110100","110100","110100","000000","000000","000000","110100","110100","110100","110100","110100","110100","111100","111100","111100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111100","111100","111100","111100","111100","110100","110100","110100","110100","110100","110100","110100","110100","110100","111100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111100","111100","111100","111100","111100","110100","110100","110100","110100","110100","110100","110100","110100","110100","111100","111100","111100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","111111","000000","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111100","111100","111100","111100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","111100","111100","111100","111100","110100","110100","110100","110100","110100","110100","110100","110100","000000","111111","111111","000000","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111100","111100","111100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","111100","111100","111100","111100","111100","110100","110100","110100","110100","000000","111111","111111","111100","000000","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111100","111100","110100","110100","110100","110100","110100","111100","110100","111100","110100","110100","110100","110100","110100","110100","110100","110100","110100","111100","111100","111100","110100","110100","110100","000000","111111","111100","111100","000000","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","111100","110100","110100","110100","110100","111100","110100","111100","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","110100","111100","110100","110100","110100","000000","111100","111100","111100","110100","000000","110100","110100","110100","000000","000000","000000","000000","000000","110100","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","110100","111100","110100","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","111100","110100","111100","110100","110100","000000","111100","111100","111100","110100","000000","110100","110100","110100","000000","000000","000000","111111","111111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","110100","110100","111100","110100","111100","110100","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","111100","110100","111100","000000","111100","111100","111100","111100","110100","000000","110100","110100","000000","111100","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","110100","111100","111100","111100","110100","110100","110100","110100","110100","110100","110100","111100","110100","111100","110100","000000","000000","000000","000000","111100","110100","110100","110100","110100","111100","110100","110100","000000","111100","111100","111100","111100","000000","000000","000000","111100","111111","111111","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","110100","111100","111100","111100","111100","110100","110100","110100","110100","110100","110100","110100","110100","111100","110100","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","111100","111100","111100","111100","111100","111100","111100","000000","111100","000000","111100","111100","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","110100","111100","111100","111100","110100","110100","110100","000000","000000","000000","110100","110100","110100","110100","110100","000000","000000","110100","110100","000000","110100","110100","110100","110100","110100","111100","111100","111100","111100","111100","111100","111100","111100","000000","111100","111111","110100","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","110100","111100","110100","110100","110100","110100","110100","000000","000000","000000","000000","110100","110100","110100","000000","000000","110100","111100","111100","110100","110100","110100","110100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111111","111111","110100","111100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","110100","111100","111100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","111100","111100","111100","111100","110100","110100","110100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111111","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","110100","111100","111100","111100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111100","111100","111100","111100","110100","110100","110100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000000","000000","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111100","111100","110100","111100","110100","110100","110100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","111100","111100","110100","111100","110100","110100","110100","110100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000000","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","110100","110100","111100","110100","110100","110100","111100","110100","110100","110100","110100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111111","111111","111111","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","111111","111111","111111","111111","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","110100","110100","111111","111111","111111","111111","111111","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","000000","000000","000000","110100","111100","110100","110100","110100","110100","110100","110100","110100","111111","111111","111111","111111","111111","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111100","111100","111100","110100","110100","110100","111100","110100","111100","110100","110100","110100","110100","110100","110100","111111","111111","111111","111111","111111","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111111","111111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","110100","110100","111100","111100","111100","111100","111100","111100","111100","110100","111100","110100","110100","110100","110100","110100","110100","111111","111111","111111","111111","111111","111111","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","110100","111100","111100","111100","110100","110100","110100","111100","111100","111100","111100","110100","110100","110100","110100","110100","110100","110100","111111","111111","111111","111111","111111","111111","111100","111100","111100","111100","111100","111100","110100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","110100","111100","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","111100","111100","111100","111100","110100","110100","110100","110100","110100","110100","111111","111111","111111","111111","111111","111111","111100","111100","111100","111100","111100","110100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","110100","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","111100","111100","111100","111100","110100","110100","110100","110100","110100","111100","111111","111111","111111","111111","111111","111100","111100","111100","111100","111100","111100","000000","000000","000000","000000","000000","111100","111100","111100","111100","111100","111100","111100","111100","111100","111100","110100","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","111100","111100","110100","110100","110100","110100","110100","110100","111111","111111","111111","111111","111111","111111","111100","111100","111100","111100","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","111100","111100","111100","110100","000000","000000","111100","111100","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","111111","111111","111111","111111","111111","111111","111111","111100","111100","111100","111100","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111100","111100","111100","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","111100","111100","110100","110100","110100","110100","110100","110100","110100","110100","111111","111111","111111","111111","111111","111111","111111","111111","111100","111100","111100","111100","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","110100","111100","111100","111100","110100","111100","110100","110100","110100","110100","110100","110100","111111","111111","111111","111111","111111","111111","111111","111111","111111","111100","111100","111100","111100","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","110100","111100","111100","111100","111100","110100","110100","110100","110100","110100","110100","110100","111111","111111","111111","111111","111111","111111","111111","111111","111100","111100","111100","111100","111100","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","110100","111100","111100","111100","110100","110100","110100","110100","110100","110100","110100","111100","111111","111111","111111","111111","111111","111111","111111","111100","111111","111100","111100","111100","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","110100","111100","110100","110100","111100","111111","110100","110100","110100","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111100","111100","111100","111100","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111100","111111","111100","111100","111100","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111100","111111","111100","111100","111100","111100","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","110100","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111100","111111","111100","111111","111100","111100","111100","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","110100","111100","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111100","111111","111100","111111","111100","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111100","111111","111100","111111","111100","111100","111100","111100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"));

constant GaradosBackString : Pokemon :=(("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","000111","000000","000000","000000","000000","000111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000000","000111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","000000","000000","000000","000000","000111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","111111","111111","111111","111111","000000","000000","000000","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000000","000000","000111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","000000","000000","000111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","000000","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000000","000000","000000","000000","111111","111111","111111","111111","000111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000000","000000","000111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","111111","111111","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","000000","000000","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","000111","000111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000000","000000","000000","000111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","000000","000000","000111","000000","000000","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000111","000000","000000","000111","000111","000111","000111","000111","000111","000111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000111","000000","111111","111111","111111","111111","000111","000111","000111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000111","000111","111111","111111","111111","111111","111111","000111","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","000111","000111","000111","000111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000111","000111","111111","000111","000111","000111","000111","000000","000000","000000","000000","000111","000111","111111","111111","111111","111111","000111","000111","000111","000111","000111","000111","000111","000000","000000","000000","000000","000000","000000","000111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000111","111111","111111","000000","000000","000000","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000111","000111","000111","000111","000111","000111","000111","000000","000000","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000000","000000","000000","000000","000111","000000","000000","000111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","111111","111111","111111","111111","000000","000000","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000111","000111","000111","000111","000111","000111","000111","000111","000000","000000","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000000","000000","000000","000111","000000","000000","000111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","000000","000111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000000","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000000","000000","000111","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","000111","000000","000000","000000","000000","000000","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000000","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000000","000111","000000","000111","000000","000111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","000000","000111","000111","000111","000000","000000","000000","000111","000111","000111","000111","000111","000111","000111","000111","000111","000000","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000000","000111","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","000000","000111","000111","000111","111000","000111","000000","000000","000000","000000","000111","000111","000111","000111","000000","000000","000000","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","111111","000000","000000","000111","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","000000","000111","000111","000111","000111","111000","111000","000111","000000","000000","000000","000000","000000","000111","000000","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000000","000111","000111","000111","000111","000111","111111","000111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","000000","000111","000111","000111","111000","111000","111000","111000","000111","000000","000000","000000","000000","000000","000000","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000000","000111","000111","000111","000111","000111","000111","111111","000000","000111","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000111","111111","111111","111111","111111","111111","111111","000000","000111","000111","000111","000111","111000","111000","111000","111000","111000","000000","000000","000111","000111","000111","000111","000000","000000","000111","000111","000111","000111","000111","000111","000111","000000","000111","000111","000111","000111","000111","000111","111111","000111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","000000","000111","000111","000111","000111","111000","111000","111000","111000","111000","000111","000000","000111","000111","000111","000111","000111","000111","000000","000111","000111","000111","000111","000000","000000","111111","000111","000111","000111","000111","000111","000111","000111","000000","000111","000111","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000111","000111","000111","000111","000111","111000","111000","111000","111000","000111","000111","000111","000000","000000","111111","111111","000111","000111","000111","000000","000000","000111","000000","111111","111111","000111","111111","000111","000111","000111","000111","000111","000111","000000","000111","000111","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","000111","111111","000000","000000","000111","000111","000111","000111","000111","000111","111000","111000","000111","000111","000111","000111","000000","111000","000000","111111","111111","111111","000111","000111","000000","000000","111111","111111","000111","111111","000111","000111","000111","000111","000111","000111","000000","000111","000111","000111","000111","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000111","111111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","111000","111000","111000","000000","111111","111111","111111","000111","000111","000000","000111","000111","111111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000000","111000","111000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000111","111111","000111","000111","000111","000111","000111","000111","000111","000111","000000","000000","000000","000111","000111","111000","111000","111000","111000","000000","111111","111111","111111","111111","000111","000111","000000","000000","000000","000000","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000000","111000","111000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000111","000111","000111","000111","000111","000000","000000","000000","111000","111000","111000","000000","000000","111000","111000","111000","000000","111111","111111","111111","111111","111111","111111","000111","000111","000000","000111","000111","000000","000111","000111","000111","000111","000111","000111","000111","000111","000111","000000","111000","111000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000111","000111","000000","000000","000000","000000","000000","111000","111000","111000","111000","111000","111000","111000","000111","000000","000000","111000","000000","111111","111111","111111","111111","111111","111111","111111","000111","000000","000000","000111","000111","000000","000111","000111","000111","000111","000111","000111","000111","000111","000111","111000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000111","111111","000111","111111","000111","000111","000111","000111","000111","111000","111000","111000","111000","111000","111000","111000","000111","000111","000111","000000","000000","111111","111111","111111","111111","111111","111111","111111","000111","000111","000000","000111","000111","000000","000111","000111","000111","000111","000111","000111","000111","000111","000111","111000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","111111","000111","111111","000111","000111","000111","000111","111000","111000","111000","111000","111000","111000","000111","000111","000111","000111","111000","000000","000000","111111","111111","111111","111111","111111","111111","111111","000111","000111","000000","000111","000000","000111","000111","000111","000111","000111","000111","000111","000111","111000","111000","000111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000111","111111","111111","111111","111111","000111","000111","000111","000111","000111","000111","111000","111000","111000","111000","111000","000111","000111","000111","111000","111000","111000","000000","000000","111111","111111","111111","111111","111111","111111","000111","000111","000000","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","111000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000111","111111","111111","111111","000111","000111","000111","000111","000111","000111","000111","111000","111000","111000","111000","111000","000111","000111","000111","111000","111000","111000","000000","000000","111111","111111","111111","000111","000111","000111","000111","000111","000111","000000","000000","000000","000111","000111","000111","000111","000111","000111","000111","111000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000111","111111","000111","111111","000111","000111","000111","000111","000111","000111","111000","111000","111000","111000","000111","000111","000111","111000","111000","111000","000000","000000","111111","111111","000111","000111","111111","111111","111111","111111","000111","000111","000000","111111","111111","000000","000111","000111","000111","000111","000111","111000","111000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","111111","000111","111111","000111","000111","000111","000111","000111","000111","000111","000111","111000","111000","000111","000111","000111","000111","111000","111000","111000","000000","111111","000111","000111","111111","111111","111111","111111","111111","111111","000111","000000","000111","000000","000000","111111","000000","000111","000111","000111","000111","111000","111000","000111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","000111","111000","111000","000000","000000","000111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000111","000111","000111","000000","111111","000000","000111","000111","000111","111000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000111","000000","000000","000000","000000","000000","000000","000000","000111","000111","000111","000111","000111","000111","000111","000111","111000","111000","111000","000000","111111","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000111","000111","000000","111111","000000","000111","000111","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000111","111111","000111","000111","000111","000111","000111","000111","000111","000000","000000","000000","000111","000111","000111","000111","000111","111000","111000","111000","000000","111111","111111","000000","111111","111111","111111","111111","111111","111111","111111","000000","000000","000111","000000","000111","000111","000000","111111","000000","000111","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000111","111111","000111","111111","000111","000111","000111","000111","111000","111000","111000","000000","000000","000000","000111","000111","111000","111000","000000","111111","111111","111111","111111","000000","111111","111111","111111","111111","111111","111111","000000","000111","000000","000111","000000","000111","000000","111111","000000","000111","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000111","111111","000111","111111","000111","000111","000111","000111","000111","111000","111000","111000","111000","000111","000111","000000","111000","111000","111000","000000","111111","111111","111111","111111","000000","111111","111111","111111","111111","111111","000000","000000","000000","000111","000000","000111","000111","000000","111111","000000","000111","000111","111000","111000","000111","000000","000000","000000","000000","000000","000000"));

constant GlurakBackString : Pokemon :=(("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000000","111111","111111","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","110100","111111","110100","110100","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","110100","111111","110100","110100","110100","111111","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000000","111111","110100","111111","110100","110100","110100","110100","110100","110100","000000","110100","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000000","000000","000000","000000","111111","111111","110100","111111","110100","110100","110100","110100","110100","110100","000000","000000","110100","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000000","111111","111111","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000000","111111","111111","111111","110100","110100","110100","110100","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000000","111111","111111","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000000","000000","000000","000000","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","110100","110100","110100","110100","110100","110100","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000101","000000","000000","000000","000000","111111","111111","111111","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","110100","110100","110100","110100","110100","000000","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","111111","111111","111111","111111","111111","111111","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000101","000000","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","111111","000101","111111","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","000000","000000","000000","110100","110100","000000","110100","110100","110100","110100","110100","110100","000000","000000","000000","111111","111111","000101","000000","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","000000","110100","110100","110100","110100","110100","000000","110100","110100","000000","111111","111111","000000","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000000","000000","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000101","000000","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","000000","111111","111111","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","111111","000000","000000","000101","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000101","111111","111111","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","000000","000000","000000","000000","000000","000000","110100","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","110100","110100","000000","000000","000000","000000","000000","000000","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111111","110100","110100","110100","110100","110100","110100","110100","110100","000000","111111","111111","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","110100","110100","110100","110100","110100","110100","110100","110100","000000","111111","111111","111111","000000","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","110100","111111","110100","110100","110100","110100","110100","110100","110100","000000","111111","111111","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111111","110100","110100","110100","110100","110100","110100","110100","110100","000101","111111","111111","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111111","110100","111111","110100","110100","110100","110100","110100","110100","110100","110100","000000","111111","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","110100","111111","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","111111","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","110100","111111","111111","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","111111","110100","110100","110100","000000","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111111","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","111111","110100","110100","110100","110100","110100","110100","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111111","111111","111111","110100","110100","110100","110100","110100","110100","110100","110100","000000","111111","000000","111111","110100","110100","110100","110100","110100","110100","110100","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","110100","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","111111","000000","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","110100","111111","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","111111","111111","110100","110100","110100","110100","000000","110100","110100","110100","110100","110100","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","110100","111111","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","111111","000000","111111","110100","111111","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","110100","111111","111111","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","111111","111111","111111","110100","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","111111","110100","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","110100","111111","110100","111111","110100","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111111","110100","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","110100","111111","110100","111111","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111111","110100","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","110100","111111","110100","111111","110100","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","111111","110100","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","110100","111111","110100","111111","110100","111111","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","110100","110100","111111","110100","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","110100","111111","110100","111111","110100","111111","110100","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","110100","111111","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","110100","110100","111111","110100","111111","110100","111111","110100","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","110100","111111","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","110100","110100","110100","111111","110100","111111","110100","111111","110100","111111","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","110100","111111","111111","110100","110100","110100","110100","110100","110100","000000","110100","110100","110100","110100","110100","111111","110100","111111","110100","111111","110100","111111","110100","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","110100","111111","111111","110100","110100","110100","110100","110100","000000","000000","110100","110100","110100","110100","110100","110100","110100","111111","110100","111111","110100","111111","110100","110100","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","110100","110100","110100","110100","110100","000000","110100","110100","110100","110100","110100","110100","111111","110100","111111","110100","111111","110100","111111","111111","111111","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","110100","110100","110100","110100","110100","110100","000000","110100","110100","110100","110100","110100","110100","111111","110100","111111","110100","111111","110100","111111","111111","111111","110100","110100","110100","000000","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","110100","000000","000000","000000","000000","000000"));

constant KokoweiBackString : Pokemon :=(("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","000000","000000","000000","111111","001000","001000","001000","001000","000000","000000","000000","001000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","111111","111111","001000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","001000","111111","001000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","001000","111111","001000","000000","000000","000000","000000","111111","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","111111","000000","000000","000000","111111","001000","111111","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","000000","111111","000000","001000","001000","001000","001000","111111","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","000000","000000","001000","001000","001000","001000","111111","001000","111111","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","000000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","001000","001000","001000","001000","000000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","111111","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","001000","001000","001000","001000","000000","001000","001000","001000","001000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","111111","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","001000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","000000","001000","000000","001000","001000","000000","000000","000000","001000","000000","001000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","001000","111111","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","000000","001000","000000","000000","001000","000000","001000","000000","001000","000000","001000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","111111","001000","001000","001000","001000","001000","000000","000000","000000","000000","001000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","000000","001000","000000","001000","000000","000000","001000","000000","001000","000000","001000","000000","000000","001000","001000","000000","000000","000000","000000","000000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","000000","001000","000000","001000","000000","000000","000000","000000","001000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","000000","000000","000000","001000","000000","000000","000000","000000","001000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","001000","000000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","001000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","001000","111111","001000","111111","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","001000","111111","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","111111","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","001000","111111","111111","001000","001000","001000","001000","001000","001000","000000","000000","001000","001000","000000","000000","000000","000000","001000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","111111","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","111111","001000","001000","000000","000000","000000","000000","000000","001000","001000","000000","000000","001000","000000","001000","000000","001000","001000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","111111","001000","111111","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","001000","001000","001000","000000","000000","000000","111111","000000","000000","001000","001000","000000","001000","001000","001000","000000","001000","000000","001000","001000","000000","000000","000000","001000","001000","001000","000000","000000","000000","000000","001000","001000","001000","111111","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","001000","001000","000000","000000","000000","000000","000000","001000","001000","001000","000000","001000","001000","001000","001000","000000","001000","001000","000000","001000","001000","000000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","001000","001000","000000","001000","001000","000000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","111000","111000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","001000","001000","001000","001000","001000","001000","000000","001000","001000","001000","001000","001000","001000","001000","000000","111000","111000","111000","111000","111000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","001000","000000","111000","111000","000000","000000","001000","001000","001000","001000","001000","000000","000000","000000","001000","001000","001000","001000","001000","001000","000000","111000","111000","111000","111111","111111","111111","111111","000000","000000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","001000","111111","111111","001000","001000","001000","001000","001000","000000","111000","111000","111000","111000","000000","001000","001000","001000","001000","001000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","000000","111000","111111","111111","111111","111111","111111","111111","000000","000000","000000","001000","001000","001000","001000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","001000","111111","001000","001000","000000","000000","111000","111000","111000","111000","111000","000000","111111","001000","001000","001000","111111","001000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","000000","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","001000","001000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","001000","111111","001000","111111","000000","000000","111111","111000","111000","111000","111000","111000","000000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","000000","111111","111111","111111","111111","001000","111111","111111","111111","000000","000000","000000","000000","001000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","001000","001000","001000","111111","001000","000000","111111","111111","000000","111111","111111","111000","111000","111000","000000","001000","111111","001000","111111","001000","001000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","000000","111111","111111","111111","000000","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","000000","111111","001000","111000","000000","111111","111111","111111","000000","111111","000000","111111","001000","111111","001000","001000","001000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","000000","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","000000","111111","111111","111111","111111","111111","111111","111111","000000","111111","000000","001000","001000","001000","001000","001000","001000","001000","000000","000000","000000","000000","000000","000000","001000","001000","001000","001000","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","000000","000000","111111","001000","111111","111111","111111","111111","111111","111111","111000","111000","000000","001000","001000","001000","001000","001000","001000","000000","000000","001000","001000","001000","000000","000000","001000","001000","001000","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","001000","001000","001000","001000","001000","001000","000000","111111","111111","111111","000000","001000","111111","111111","111111","111111","111111","111111","000000","001000","001000","001000","001000","001000","001000","000000","001000","001000","111000","001000","111000","001000","000000","001000","001000","000000","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","001000","001000","001000","001000","001000","000000","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","111111","111000","000000","001000","001000","001000","001000","001000","001000","000000","111000","001000","111000","001000","001000","001000","000000","001000","000000","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","001000","001000","001000","001000","000000","000000","000000","111111","111111","111111","111111","001000","000000","000000","000000","000000","111111","111000","000000","001000","001000","001000","001000","001000","001000","000000","001000","111000","001000","111000","001000","111000","111000","000000","111000","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","001000","001000","001000","001000","000000","000000","001000","111111","111111","111111","111111","111111","111111","000000","000000","111111","111000","111000","111000","000000","001000","001000","001000","001000","001000","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","001000","001000","001000","001000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111000","111000","111000","000000","001000","001000","001000","001000","001000","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","001000","001000","001000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111000","111000","111000","111000","111000","000000","001000","001000","001000","001000","001000","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","001000","001000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111000","111000","111000","111000","111000","000000","000000","000000","001000","001000","001000","001000","000000","111000","111000","111000","111000","111000","111000","111000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","001000","001000","000000","000000","000000","000000","000000","000000","000000","001000","000000","111000","111000","111000","111000","111000","000000","000000","111000","111000","000000","000000","001000","001000","001000","000000","111000","111000","111000","111000","111000","111000","111000","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","111000","111000","111000","111000","000000","000000","001000","001000","001000","000000","111000","111000","111000","111000","000000","000000","111000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111000","000000","000000","000000","111000","111000","111000","111000","111000","000000","001000","001000","000000","111000","000000","000000","000000","111000","111000","111111","111000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111000","111111","111000","111000","111000","001000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","111000","111000","111000","111111","111000","111111","111000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","111111","111000","111111","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111111","111000","111111","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"));

constant MagmarBackString : Pokemon :=(("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","000000","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","000000","000000","100101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111000","111111","111000","111111","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","111111","000000","111111","111111","111111","111111","000000","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","111111","111000","111111","111000","111111","111000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111000","111111","111000","111111","111000","111111","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111000","111111","111000","000000","000000","000000","000000","000000","000000","100101","000000","111000","111000","111111","111000","111111","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111000","111111","111000","111111","111000","000000","000000","000000","000000","000000","000000","000000","111000","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","111111","111000","111111","111000","000000","000000","000000","000000","000000","000000","100101","111000","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","111111","111000","111111","000000","000000","000000","000000","000000","000000","000000","111000","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","111000","111000","111000","000000","000000","111000","111000","000000","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","111000","111000","111000","111000","111000","111000","111000","100101","100101","100101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","111000","111000","111000","111000","111000","111000","100101","111000","100101","100101","100101","100101","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","111000","111000","111000","111000","111000","111000","100101","111000","100101","111000","100101","100101","100101","100101","111000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","100101","111111","111111","111000","111000","111000","111000","111000","111000","100101","111000","100101","100101","100101","100101","111000","100101","111000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","111000","111000","000000","111000","111000","111000","111000","111000","111111","111111","111000","111111","111000","111000","111000","111000","100101","111000","100101","100101","100101","100101","100101","100101","111000","100101","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","111000","111000","111000","111000","111111","111111","111000","111111","111000","111000","111000","111000","111000","111000","100101","100101","100101","100101","100101","100101","111000","100101","111000","100101","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","111000","111000","111000","111000","111111","111000","111111","111000","111111","111000","111000","111000","111000","111000","100101","100101","100101","100101","100101","100101","100101","111000","100101","111000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","111000","111000","111000","000000","000000","000000","100101","000000","000000","000000","000000","000000","100101","111000","111000","111000","111000","111000","111000","111000","111111","111000","111111","111000","111000","111000","111000","111000","111000","111000","100101","100101","100101","100101","100101","100101","100101","111000","100101","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","100101","100101","100101","100101","111000","111000","000000","000000","000000","100101","000000","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","100101","100101","100101","100101","100101","100101","100101","100101","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","100101","100101","100101","100101","100101","100101","100101","111000","111000","000000","000000","000000","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","100101","000000","100101","100101","100101","100101","100101","100101","100101","100101","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","000000","000000","000000","111000","111000","111000","111000","111000","111000","111000","100101","111000","100101","100101","100101","000000","000000","111111","111111","100101","100101","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","000000","111000","100101","111000","100101","111000","100101","111000","100101","100101","100101","100101","100101","100101","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","000000","100101","111000","100101","111000","100101","111000","100101","111000","100101","100101","100101","100101","100101","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","000000","100101","100101","111000","100101","111000","100101","100101","100101","100101","100101","100101","100101","100101","000000","111111","000000","111000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","100101","100101","100101","100101","100101","100101","000000","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","000000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","111000","111000","000000","100101","100101","100101","100101","100101","100101","000000","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","000000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","111111","111111","111111","111000","111000","000000","000000","100101","100101","100101","100101","000000","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","000000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","100101","000000","000000","000000","000000","000000","111000","111111","111111","111111","111111","111000","111000","111000","000000","000000","000000","100101","000000","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","000000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","100101","111000","111000","111000","111000","100101","100101","000000","000000","000000","000000","000000","000000","000000","111000","000000","000000","000000","000000","000000","000000","100101","100101","100101","100101","100101","000000","000000","000000","000000","000000","000000","100101","100101","000000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","000000","000000","000000","000000","000000","000000","100101","100101","100101","100101","000000","000000","111000","111000","111000","111000","111000","111000","000000","000000","111000","111000","111000","100101","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","000000","000000","000000","000000","000000","100101","000000","111000","111000","111111","111111","111111","111000","111000","111000","111000","111000","000000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","000000","000000","000000","000000","000000","000000","111000","111000","111111","111111","111111","111111","111111","111000","111000","111000","111000","111000","000000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","100101","100101","100101","100101","100101","100101","100101","100101","000000","000000","000000","000000","000000","000000","111000","111000","111111","111111","111111","111111","111111","111111","111000","111000","111000","111000","111000","111000","000000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","100101","100101","100101","100101","100101","100101","000000","000000","000000","000000","000000","000000","111000","111000","111111","111111","111111","111111","111111","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","111000","000000","000000","100101","100101","100101","100101","000000","000000","000000","000000","000000","000000","111000","111000","111000","111000","111111","111111","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","111000","111000","111000","000000","000000","100101","100101","000000","100101","100101","000000","000000","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","100101","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111000","111000","111000","000000","100101","000000","000000","100101","100101","100101","100101","100101","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","100101","111000","111000","111000","111000","100101","100101","100101","100101","000000","000000","000000","000000","000000","000000","000000","000000","100101","100101","100101","100101","100101","100101","100101","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","111000","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","000000","100101","100101","100101","100101","100101","100101","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","000000","100101","100101","100101","100101","100101","100101","100101","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","100101","000000","100101","100101","100101","100101","100101","100101","100101","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","100101","100101","100101","100101","100101","100101","000000","100101","100101","100101","100101","111000","100101","111000","100101","100101","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","100101","000000","100101","100101","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","100101","100101","100101","100101","000000","100101","100101","100101","111000","100101","111000","100101","100101","100101","100101","000000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","100101","100101","000000","100101","100101","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","100101","100101","000000","100101","100101","111000","100101","111000","100101","111000","100101","100101","100101","100101","000000","000000","111000","111000","111000","111000","111000","111000","000000","000000","100101","000000","100101","100101","000000","100101","100101","000000","000000","000000","000000","000000","000000","000000"));

constant SarzeniaBackString : Pokemon :=(("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","011100","011100","011100","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","000000","000000","111111","111111","111111","011100","011100","011100","000000","000000","000000","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","011100","011100","011100","011100","011100","011100","000000","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","011100","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","011100","011100","011100","011100","011100","011100","000000","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","000000","000000","000000","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","011100","011100","111111","011100","111111","011100","000000","000000","011100","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","111111","111111","111111","111111","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","011100","000000","011100","111111","011100","111111","011100","111111","000000","011100","000000","011100","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","011100","111111","011100","111111","011100","111111","000000","011100","000000","011100","000000","011100","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","011100","000000","111111","011100","111111","011100","111111","011100","000000","000000","011100","000000","011100","000000","011100","000000","011100","011100","011100","000000","000000","000000","000000","000000","000000","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","111111","011100","000000","011100","111111","011100","111111","011100","000000","000000","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","110110","110110","110110","110110","111111","111111","000000","000000","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","111111","111111","011100","000000","111111","011100","111111","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","110110","110110","110110","110110","110110","110110","110110","110110","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","111111","111111","000000","011100","011100","111111","011100","011100","000000","000000","000000","000000","000000","000000","000000","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","111111","011100","000000","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","111111","110110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","011100","000000","111111","011100","000000","011100","011100","011100","011100","011100","000000","000000","000000","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","111111","110110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","011100","111111","000000","111111","011100","011100","011100","011100","011100","011100","011100","000000","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","110110","000000","000000","000000","000000","000000","000000","000000","110110","110110","110110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","011100","011100","000000","111111","011100","000000","011100","011100","011100","011100","000000","110110","110110","110110","110110","110110","110110","110110","110110","110110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","000000","110110","110110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","011100","011100","000000","111111","011100","011100","011100","011100","011100","011100","000000","110110","110110","110110","110110","110110","110110","110110","000000","000000","000000","000000","000000","110110","011100","011100","011100","110110","000000","000000","111111","000000","110110","110110","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","011100","011100","000000","111111","011100","000000","011100","011100","011100","000000","110110","110110","110110","110110","110110","110110","000000","000000","000000","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","011100","000000","111111","011100","011100","011100","011100","011100","000000","110110","110110","110110","110110","110110","000000","000000","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","011100","000000","111111","011100","000000","011100","011100","000000","110110","110110","110110","110110","000000","000000","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","111111","111111","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","011100","000000","111111","011100","000000","011100","000000","110110","110110","110110","110110","000000","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","111111","111111","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","000000","110110","110110","110110","110110","000000","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","111111","111111","111111","011100","000000","111111","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","000000","110110","110110","110110","000000","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","111111","111111","011100","000000","110110","110110","000000","000000","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","011100","000000","110110","110110","000000","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","000000","110110","110110","000000","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","111111","111111","111111","111111","111111","111111","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","111111","111111","000000","000000","000000","000000","000000","011100","011100","111111","011100","111111","011100","111111","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","011100","000000","000000","000000","000000","000000","111111","011100","111111","011100","111111","011100","111111","011100","011100","011100","011100","011100","011100","011100","011100","011100","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","000000","000000","000000","000000","000000","000000","111111","011100","111111","011100","111111","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","111111","111111","111111","111111","111111","111111","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","111111","111111","011100","000000","000000","000000","000000","000000","011100","111111","011100","111111","011100","111111","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","111111","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","000000","000000","000000","000000","000000","000000","011100","111111","011100","111111","011100","111111","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","111111","111111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","011100","000000","000000","000000","000000","000000","111111","011100","111111","011100","111111","011100","011100","011100","011100","011100","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","000000","000000","000000","000000","000000","000000","111111","011100","111111","011100","111111","011100","111111","011100","111111","011100","011100","000000","000000","000000","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","011100","000000","011100","011100","011100","000000","011100","111111","011100","111111","011100","111111","011100","111111","011100","000000","000000","011100","011100","011100","011100","000000","000000","111111","111111","111111","111111","111111","000000","011100","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","011100","000000","011100","011100","000000","111111","011100","111111","011100","111111","011100","111111","011100","000000","011100","011100","011100","011100","011100","111111","111111","111111","000000","000000","111111","111111","111111","111111","111111","000000","011100","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","011100","000000","011100","011100","000000","111111","011100","111111","011100","111111","011100","000000","011100","011100","011100","011100","111111","111111","111111","111111","111111","111111","011100","000000","011100","011100","011100","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","011100","011100","000000","011100","011100","011100","000000","011100","000000","011100","111111","011100","111111","011100","000000","011100","011100","111111","111111","111111","111111","111111","111111","011100","011100","011100","011100","011100","000000","011100","011100","011100","011100","011100","011100","000000","000000","000000","000000","000000","000000","000000"));

constant TurtokBackString : Pokemon :=(("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","000000","111111","111111","111111","010111","010111","000000","000000","010111","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","010111","010111","010111","000000","000000","010111","111111","111111","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","000000","000000","000000","010111","111111","111111","111111","111111","111111","111111","111111","010111","111111","010111","010111","010111","010111","000000","000000","010111","010111","010111","010111","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","111111","111111","010111","010111","010111","010111","111111","111111","111111","111111","111111","111111","010111","111111","010111","010111","010111","010111","010111","010111","010111","000000","000000","010111","010111","010111","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","111111","010111","010111","010111","010111","111111","111111","111111","111111","111111","111111","010111","111111","010111","010111","010111","010111","010111","010111","010111","111111","111111","010111","010111","010111","010111","010111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","010111","010111","010111","010111","111111","111111","111111","010111","111111","010111","111111","010111","010111","010111","000000","000000","000000","000000","111111","111111","111111","010111","010111","000000","010111","010111","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","010111","010111","010111","010111","010111","111111","010111","111111","010111","111111","010111","010111","010111","010111","010111","010111","010111","010111","000000","111111","010111","010111","000000","000000","000000","010111","010111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","010111","010111","010111","010111","010111","111111","010111","010111","010111","010111","010111","010111","010111","111111","111111","010111","010111","010111","010111","000000","000000","000000","000000","010111","010111","010111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","111111","111111","111000","010111","000000","000000","010111","000000","111111","111111","000000","010111","010111","010111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","111000","111000","010111","000000","000000","000000","010111","000000","111111","111111","000000","010111","010111","010111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","010111","000000","111111","111111","111111","111111","000000","010111","000000","000000","000000","000000","000000","000000","000000","000000","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","000000","000000","010111","010111","010111","111111","000000","010111","010111","010111","010111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","010111","111111","111111","111111","111000","010111","010111","111111","111111","010111","000000","000000","000000","000000","000000","000000","000000","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","111111","000000","010111","010111","010111","010111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111000","010111","010111","010111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","000000","010111","010111","010111","010111","000000","010111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","010111","111111","111111","111111","111111","111000","010111","010111","111111","010111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","000000","000000","000000","010111","010111","010111","010111","010111","010111","010111","010111","010111","010111","000000","010111","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111000","010111","010111","010111","111111","010111","000000","000000","000000","000000","010111","000000","111111","111111","111111","111111","000000","000000","000000","010111","010111","010111","010111","010111","010111","000000","111111","111111","111111","000000","000000","010111","010111","010111","010111","010111","010111","010111","000000","111111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111000","010111","010111","111111","010111","111111","000000","000000","000000","000000","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","010111","010111","010111","000000","111111","010111","000000","000000","111111","111111","000000","000000","010111","010111","010111","010111","000000","111000","111111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111000","010111","010111","010111","111111","010111","000000","000000","010111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","010111","010111","000000","111111","111111","000000","000000","000000","000000","111111","111111","000000","010111","010111","000000","111000","111000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","111111","111111","111111","111000","010111","010111","111111","010111","111111","000000","000000","000000","000000","000000","000000","010111","111111","111111","111111","111111","111111","111111","111111","111111","111111","000000","000000","111111","111111","111111","111111","000000","000000","000000","000000","111111","111111","000000","010111","000000","111000","111000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","000000","111111","010111","000000","000000","000000","010111","010111","010111","111111","010111","000000","111000","111111","111000","111111","111000","111000","000000","000000","010111","111111","111111","111111","111111","111111","111000","111111","000000","111111","111111","111111","111111","111111","000000","000000","000000","000000","111111","000000","000000","111000","111000","111000","010111","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","010111","000000","111111","111000","111000","111000","000000","000000","000000","000000","111000","111000","111111","111111","111111","111000","111000","111000","111000","111000","111000","000000","000000","111111","111111","111000","111111","000000","111111","111111","111111","111111","111111","111111","111111","010111","000000","000000","000000","111111","000000","111000","111000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","010111","111111","111111","111111","111000","111000","111000","111000","000000","111000","111000","111111","111111","111111","111111","111000","111111","111000","111000","111000","111000","111000","111000","111000","000000","000000","111111","111000","000000","111111","111111","111111","111111","111111","111000","010111","111111","111111","010111","010111","111111","000000","111000","111000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","111111","111111","111000","111000","111000","111000","000000","111000","111000","111111","111111","111111","111111","111000","111111","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","000000","111111","111111","111111","111111","111111","111111","010111","010111","010111","111111","111111","111111","111111","000000","111000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","010111","111111","111111","111111","111000","111000","111000","000000","111000","111000","111111","111111","111111","111111","111000","111111","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","111111","111111","111111","111111","111111","111000","010111","010111","111111","010111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","111111","111111","111111","111000","111000","000000","111000","111000","000000","000000","000000","000000","010111","111111","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","111111","111111","111111","111111","111111","111111","010111","010111","111111","010111","111111","111111","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","111111","111111","111000","111000","000000","111000","000000","000000","111000","111111","111111","111111","000000","000000","000000","000000","010111","111000","111000","111000","111000","111000","111000","000000","000000","000000","000000","111111","111111","111111","111111","111111","111000","010111","111111","010111","111111","010111","111111","000000","000000","010111","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","111111","111111","111000","111000","000000","000000","111000","111111","111111","111111","111111","111111","111000","111111","111000","111000","000000","000000","010111","010111","111000","000000","000000","111111","111111","111111","000000","000000","111111","111111","111111","111111","010111","010111","010111","111111","010111","111111","111111","000000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","111111","111111","111000","000000","111000","111111","111111","111111","111111","111111","111111","111000","111111","111000","111000","111000","111000","111000","000000","000000","000000","010111","111111","111111","111111","111111","111111","000000","000000","111111","111111","111000","010111","010111","111111","010111","111111","111111","000000","111111","111000","111111","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","111111","111111","000000","111000","111000","111111","111111","111111","111111","111111","111000","111111","111000","111000","111000","111000","111000","111000","111000","000000","000000","111111","111111","111111","111111","111111","111111","111111","000000","000000","111111","010111","010111","111111","010111","111111","010111","111111","000000","111000","111111","111000","111111","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","010111","111111","111111","000000","111000","111111","111111","111111","111111","111111","111000","111111","111000","111111","111000","111000","111000","111000","111000","111000","111000","000000","111111","111111","111000","111000","111000","111111","111111","111111","010111","000000","000000","010111","010111","111111","010111","111111","000000","000000","111111","111000","111111","111000","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","010111","000000","111000","111000","111111","111111","111111","111111","111000","111111","111000","111111","111000","111000","111000","111000","111000","111000","111000","010111","111111","111111","111000","111000","111000","111000","111000","111000","111111","111111","111111","010111","000000","000000","111111","111111","000000","000000","000000","000000","000000","111000","111111","111111","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","010111","000000","111000","111000","111111","111111","111111","111000","111111","111000","111111","111000","111000","111000","111000","111000","111000","111000","111000","000000","111111","111111","111000","111000","111000","111000","111000","111000","111000","111000","111111","111111","111000","010111","000000","000000","000000","000000","010111","010111","010111","000000","000000","111111","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","010111","000000","111000","111111","111111","111111","111000","111111","111000","111111","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","111111","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","010111","000000","010111","111111","111111","010111","010111","010111","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","111000","111000","111111","111111","111000","111111","111000","111111","111000","111111","111000","111000","111000","111000","111000","111000","111000","010111","111111","111111","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","111111","111111","010111","010111","010111","000000","000000","000000","000000","000000","000000","000000","000000"),
("000000","000000","000000","000000","000000","000000","111000","111000","111111","111111","111111","111000","111111","111000","111111","111000","111000","111000","111000","111000","111000","111000","111000","000000","111111","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","111000","000000","010111","010111","010111","010111","010111","010111","000000","000000","000000","000000","000000","000000","000000"));


signal limit: integer;
signal Hp1 : integer;
signal Hp2 : integer;

begin

Hp1 <= 2 * to_integer(unsigned(t1p1(8 downto 4)));
Hp2 <= 2 * to_integer(unsigned(t2p1(8 downto 4)));

process (display)

variable rot : integer := to_integer(unsigned(sschaden)) + to_integer(unsigned(sschaden));
variable pixelX : integer := to_integer(unsigned(pixel_X));
variable pixelY : integer := to_integer(unsigned(pixel_Y));

begin


if(display ='1' and rising_edge(Halfclock)) then
    
    --resets the colors
     rin <= "0000";
     gin <= "0000";
     bin <= "0000";
    
    --The Main Menu
    if (menu = "000")then  
        
        if(pixel_x > 259  and pixel_x < 541  and pixel_y > 50 and pixel_y < 210) then --Pokemon yaz�s�
    
            rin(3 downto 2) <= PokemonString (pixelY - 51, pixelX - 260) (5 downto 4);
            gin(3 downto 2) <= PokemonString (pixelY - 51, pixelX - 260) (3 downto 2);
            bin(3 downto 2) <= PokemonString (pixelY - 51, pixelX - 260) (1 downto 0);
        elsif(pixel_x > 160  and pixel_x < 292  and pixel_y > 400 and pixel_y < 427) then --singleplayer yaz�s�
        
            if(singleplayerstring(PixelY- 401,pixelX-161) = '0') then
            rin <= "0000";
            gin <= "0000";
            bin <= "0000";
            else
            rin <= "1111";
            gin <= "1111";
            bin <= "0000";
            end if;
           
        elsif(pixel_x > 550  and pixel_x < 675  and pixel_y > 400 and pixel_y < 427) then --multiplayer yaz�s�
            
            if(multiplayerstring(PixelY- 401,pixelX-551) = '0') then
            rin <= "0000";
            gin <= "0000";
            bin <= "0000";
            else
            rin <= "1111";
            gin <= "1111";
            bin <= "0000";
            end if;
            
         else 
         
            rin <= "0000";
            gin <= "0000";
            bin <= "0000";    
        end if; -- the menu ends
            
     --Single or Multi PokemonChoice Screen
     elsif (menu = "001" or menu = "010" )then       
        
        --HP
        if (pixelY > 176 and pixelY < 233 and pixelX > 20 and pixelX < 83) then             
            rin(3 downto 2) <= HpString (pixelY - 176, pixelX - 20) (5 downto 4);
            gin(3 downto 2) <= HpString (pixelY - 176, pixelX - 20) (3 downto 2);
            bin(3 downto 2) <= HpString (pixelY - 176, pixelX - 20) (1 downto 0);
        
        limit <= to_integer(unsigned(PokemonStats(19 downto 15)));    
        elsif (pixelY > 203 and pixelY < 208 and pixelX > 110 and pixelX < 110 + 2*limit) then
            rin <= "1111";
            gin <= "1111";
            bin <= "1111";
        
        --AT
        elsif (pixelY > 243 and pixelY < 295 and pixelX > 20 and pixelX < 91) then
            rin(3 downto 2) <= AtString (pixelY - 243, pixelX - 20) (5 downto 4);
            gin(3 downto 2) <= AtString (pixelY - 243, pixelX - 20) (3 downto 2);
            bin(3 downto 2) <= AtString (pixelY - 243, pixelX - 20) (1 downto 0);
        
        limit <= to_integer(unsigned(PokemonStats(14 downto 10)));    
        elsif (pixelY > 268 and pixelY < 273 and pixelX > 110 and pixelX < 110 + 2*limit) then
            rin <= "1111";
            gin <= "1111";
            bin <= "1111";
                            
        --DEF
        elsif (pixelY > 305 and pixelY < 350 and pixelX > 20 and pixelX < 102) then
            rin(3 downto 2) <= DefString (pixelY - 305, pixelX - 20) (5 downto 4);
            gin(3 downto 2) <= DefString (pixelY - 305, pixelX - 20) (3 downto 2);
            bin(3 downto 2) <= DefString (pixelY - 305, pixelX - 20) (1 downto 0);
        
        limit <= to_integer(unsigned(PokemonStats(9 downto 5)));    
        elsif (pixelY > 326 and pixelY < 331 and pixelX > 110 and pixelX < 110 + 2*limit) then
            rin <= "1111";
            gin <= "1111";
            bin <= "1111";
                    
        --SP
        elsif (pixelY > 360 and pixelY < 415 and pixelX > 20 and pixelX < 83) then
            rin(3 downto 2) <= SpString (pixelY - 360, pixelX - 20) (5 downto 4);
            gin(3 downto 2) <= SpString (pixelY - 360, pixelX - 20) (3 downto 2);
            bin(3 downto 2) <= SpString (pixelY - 360, pixelX - 20) (1 downto 0);
        
        limit <= to_integer(unsigned(PokemonStats(4 downto 0)));    
        elsif (pixelY > 387 and pixelY < 392 and pixelX > 110 and pixelX < 110 + 2*limit) then
            rin <= "1111";
            gin <= "1111";
            bin <= "1111";
        
        --Pokemon Pictures 
        elsif (pixelY > 202 and pixelY < 258) then
        
            if (pixelX > 260  and pixelX < 316) then
            
                rin(3 downto 2) <=  AustossFrontString(pixelY - 140, pixelX - 261) (5 downto 4);
                gin(3 downto 2) <=  AustossFrontString(pixelY - 140, pixelX - 261) (3 downto 2);
                bin(3 downto 2) <=  AustossFrontString(pixelY - 140, pixelX - 261) (1 downto 0);
            
            elsif(pixelX > 372 and pixelX < 428) then
            
                rin(3 downto 2) <=  GaradosFrontString(pixelY - 140, pixelX - 373) (5 downto 4);
                gin(3 downto 2) <=  GaradosFrontString(pixelY - 140, pixelX - 373) (3 downto 2);
                bin(3 downto 2) <=  GaradosFrontString(pixelY - 140, pixelX - 373) (1 downto 0);
            
            elsif (pixelX > 484  and pixelX < 540) then
            
                rin(3 downto 2) <=  TurtokFrontString(pixelY - 140, pixelX - 485) (5 downto 4);
                gin(3 downto 2) <=  TurtokFrontString(pixelY - 140, pixelX - 485) (3 downto 2);
                bin(3 downto 2) <=  TurtokFrontString(pixelY - 140, pixelX - 485) (1 downto 0);
            
            else
            
                rin <= "0000";
                gin <= "0000";
                bin <= "0000";
            
            end if;  
        
        elsif(pixelY > 272 and pixelY < 328) then 
        
            if (pixelX > 260 and pixelX < 316) then
                    
                rin(3 downto 2) <=  BisaflorFrontString(pixelY - 210, pixelX - 261) (5 downto 4);
                gin(3 downto 2) <=  BisaflorFrontString(pixelY - 210, pixelX - 261) (3 downto 2);
                bin(3 downto 2) <=  BisaflorFrontString(pixelY - 210, pixelX - 261) (1 downto 0);
            
            elsif(pixelX > 372  and pixelX < 428) then
            
                rin(3 downto 2) <=  KokoweiFrontString(pixelY - 210, pixelX - 373) (5 downto 4);
                gin(3 downto 2) <=  KokoweiFrontString(pixelY - 210, pixelX - 373) (3 downto 2);
                bin(3 downto 2) <=  KokoweiFrontString(pixelY - 210, pixelX - 373) (1 downto 0);
            
            elsif (pixelX > 484  and pixelX < 540) then
            
                rin(3 downto 2) <=  SarzeniaFrontString(pixelY - 210, pixelX - 485) (5 downto 4);
                gin(3 downto 2) <=  SarzeniaFrontString(pixelY - 210, pixelX - 485) (3 downto 2);
                bin(3 downto 2) <=  SarzeniaFrontString(pixelY - 210, pixelX - 485) (1 downto 0);
            
            else
            
                rin <= "0000";
                gin <= "0000";
                bin <= "0000";
            
            end if;
        
        elsif(pixelY > 342 and pixelY < 398) then
        
            if (pixelX > 260  and pixelX < 316) then
                    
                rin(3 downto 2) <=  GlurakFrontString(pixelY - 280, pixelX - 261) (5 downto 4);
                gin(3 downto 2) <=  GlurakFrontString(pixelY - 280, pixelX - 261) (3 downto 2);
                bin(3 downto 2) <=  GlurakFrontString(pixelY - 280, pixelX - 261) (1 downto 0);
            
            elsif(pixelX > 372  and pixelX < 428) then
            
                rin(3 downto 2) <=  MagmarFrontString(pixelY - 280, pixelX - 373) (5 downto 4);
                gin(3 downto 2) <=  MagmarFrontString(pixelY - 280, pixelX - 373) (3 downto 2);
                bin(3 downto 2) <=  MagmarFrontString(pixelY - 280, pixelX - 373) (1 downto 0);
            
            elsif (pixelX > 484  and pixelX < 540) then
            
                rin(3 downto 2) <=  GallopaFrontString(pixelY - 280, pixelX - 485) (5 downto 4);
                gin(3 downto 2) <=  GallopaFrontString(pixelY - 280, pixelX - 485) (3 downto 2);
                bin(3 downto 2) <=  GallopaFrontString(pixelY - 280, pixelX - 485) (1 downto 0);
            
            else
            
                rin <= "0000";
                gin <= "0000";
                bin <= "0000";
            
            end if;
        
        end if;
        --Pokemon Chooser Frame       
        if((pixelY > 194  and pixelY < 198) or (pixelY > 261 and pixelY < 265)) then
            
            if((((pixelX > 251 and pixelX < 255) or (pixelX > 321 and pixelX < 325)) and pokemonchooser = 0) or (pokemonFramer(0) = '1' and ((pixelX > 251 and pixelX < 255) or (pixelX > 321 and pixelX < 325)))) then
            rin <= "1111";
                            gin <= "1111";
                            bin <= "1111";
            end if;
            if((((pixelX > 363 and pixelX < 367) or (pixelX > 433 and pixelX < 437)) and pokemonchooser = 1) or (pokemonFramer(1) = '1' and ((pixelX > 363 and pixelX < 367) or (pixelX > 433 and pixelX < 437)))) then
            rin <= "1111";
                                            gin <= "1111";
                                            bin <= "1111";
            end if;
            if((((pixelX > 475 and pixelX < 479) or (pixelX > 545 and pixelX < 549)) and pokemonchooser = 2) or (((pixelX > 475 and pixelX < 479) or (pixelX > 545 and pixelX < 549)) and pokemonFramer(2) = '1')) then
            rin <= "1111";
                                            gin <= "1111";
                                            bin <= "1111";       
            end if;
            
         end if;

        if((pixelY > 275 and pixelY < 279) or (pixelY > 331 and pixelY < 335)) then
            
            if((((pixelX > 251 and pixelX < 255) or (pixelX > 321 and pixelX < 325)) and pokemonchooser = 3) or (pokemonFramer(3) = '1' and ((pixelX > 251 and pixelX < 255) or (pixelX > 321 and pixelX < 325)))) then
            rin <= "1111";
                                            gin <= "1111";
                                            bin <= "1111";
            end if;            
            if((((pixelX > 363 and pixelX < 367) or (pixelX > 433 and pixelX < 437)) and pokemonchooser = 4) or (pokemonFramer(4) = '1' and ((pixelX > 363 and pixelX < 367) or (pixelX > 433 and pixelX < 437)))) then
            rin <= "1111";
                                            gin <= "1111";
                                            bin <= "1111";
            end if;
            if((((pixelX > 475 and pixelX < 479) or (pixelX > 545 and pixelX < 549)) and pokemonchooser = 5) or (((pixelX > 475 and pixelX < 479) or (pixelX > 545 and pixelX < 549)) and pokemonFramer(5) = '1')) then
            rin <= "1111";
                                            gin <= "1111";
                                            bin <= "1111";
            end if;
            
        end if;
        
        if((pixelY > 341 and pixelY < 345) or (pixelY > 401 and pixelY < 405)) then
        
           if((((pixelX > 251 and pixelX < 255) or (pixelX > 321 and pixelX < 325)) and pokemonchooser = 6) or (pokemonFramer(6) = '1' and ((pixelX > 251 and pixelX < 255) or (pixelX > 321 and pixelX < 325)))) then
           rin <= "1111";
                                           gin <= "1111";
                                           bin <= "1111";
           end if;             
           if((((pixelX > 363 and pixelX < 367) or (pixelX > 433 and pixelX < 437)) and pokemonchooser = 7) or (pokemonFramer(7) = '1' and ((pixelX > 363 and pixelX < 367) or (pixelX > 433 and pixelX < 437)))) then
           rin <= "1111";
                                           gin <= "1111";
                                           bin <= "1111";
           end if; 
           if((((pixelX > 475 and pixelX < 479) or (pixelX > 545 and pixelX < 549)) and pokemonchooser = 8) or (((pixelX > 475 and pixelX < 479) or (pixelX > 545 and pixelX < 549)) and pokemonFramer(8) = '1')) then
           rin <= "1111";
                                           gin <= "1111";
                                           bin <= "1111";
           end if;
            
         end if;
            
           
            --Choose
            if(pixelx > 288 and pixelx < 400 and pixely >100 and pixely <138) then
                if(Choosestring(pixely-101, pixelx-289) = '0')then
                rin <= "0000";
                gin <= "0000";
                bin <= "0000";
                else
                rin <= "1111";
                gin <= "1111";
                bin <= "1111";
                end if;
                
            --Team
            elsif(pixelx > 403 and pixelx < 491 and pixely >100 and pixely <134) then
                if(teamstring(pixely-101, pixelx-404) = '0')then
                rin <= "0000";
                gin <= "0000";
                bin <= "0000";
                else
                rin <= "1111";
                gin <= "1111";
                bin <= "1111";
                end if;
            --1 or 2
            elsif(pixely >100 and pixely <134) then
                if(Pokemonnumbers < 2 or ssingle = '1') then
                    if(pixelx > 493 and pixelx < 509) then
                        if(onestring(pixely-101, pixelx-494) = '0')then
                        rin <= "0000";
                        gin <= "0000";
                        bin <= "0000";
                        else
                        rin <= "1111";
                        gin <= "1111";
                        bin <= "1111";
                        end if;
                    end if;
                 else
                    if(pixelx > 493 and pixelx < 515) then
                         if(twostring(pixely-101, pixelx-494) = '0')then
                         rin <= "0000";
                         gin <= "0000";
                         bin <= "0000";
                         else
                         rin <= "1111";
                         gin <= "1111";
                         bin <= "1111";
                         end if;
                     end if;
                  end if;
            end if;
            
     --Single or Multi Fight
     elsif (menu = "011" or menu = "100") then
     
          --White Lines
          if((pixelY > 400 and pixelY < 405 and PixelX > 150 and PixelX < 650)  or (pixelY > 500 and pixelY < 505 and PixelX > 150 and PixelX < 650)) then
              rin <= "1111";
              gin <= "1111";
              bin <= "1111";
              
          --HP1    
          elsif(pixelY > 283 and pixelY < 340 and PixelX > 200 and PixelX < 266 and PAliveStatus(0) = '1') then
            rin(3 downto 2) <= HpString (pixelY - 284, pixelX - 201) (5 downto 4);
            gin(3 downto 2) <= HpString (pixelY - 284, pixelX - 201) (3 downto 2);
            bin(3 downto 2) <= HpString (pixelY - 284, pixelX - 201) (1 downto 0);
            
             
          elsif (pixelY > 309 and pixelY < 313 and pixelX > 270 and pixelX < 270 + hp1) then
            rin <= "1111";
            gin <= "1111";
            bin <= "1111";
          
          --HP2
          elsif(pixelY > 153 and pixelY < 210 and PixelX > 470 and PixelX < 536 and PAliveStatus(2) = '1') then
            rin(3 downto 2) <= HpString (pixelY - 154, pixelX - 471) (5 downto 4);
            gin(3 downto 2) <= HpString (pixelY - 154, pixelX - 471) (3 downto 2);
            bin(3 downto 2) <= HpString (pixelY - 154, pixelX - 471) (1 downto 0);
          
          elsif (pixelY > 179 and pixelY < 183 and pixelX > 540 and pixelX < 540 + hp2) then
            rin <= "1111";
            gin <= "1111";
            bin <= "1111";
      
          
          --T1P1
          elsif(pixelY > 344 and pixelY < 401 and PixelX > 230 and PixelX < 286 and PAliveStatus(0) = '1') then
             if(t1p1(3 downto 0) = "0000") then
                          rin(3 downto 2) <=  AustossbackString(pixelY - 345, pixelX - 231) (5 downto 4);
                          gin(3 downto 2) <=  AustossbackString(pixelY - 345, pixelX - 231) (3 downto 2);
                          bin(3 downto 2) <=  AustossbackString(pixelY - 345, pixelX - 231) (1 downto 0); 
              elsif(t1p1(3 downto 0) = "0001") then
                           rin(3 downto 2) <=  GaradosbackString(pixelY - 345, pixelX - 231) (5 downto 4);
                           gin(3 downto 2) <=  GaradosbackString(pixelY - 345, pixelX - 231) (3 downto 2);
                           bin(3 downto 2) <=  GaradosbackString(pixelY - 345, pixelX - 231) (1 downto 0);
              elsif(t1p1(3 downto 0) = "0010") then 
                           rin(3 downto 2) <=  TurtokbackString(pixelY - 345, pixelX - 231) (5 downto 4);
                           gin(3 downto 2) <=  TurtokbackString(pixelY - 345, pixelX - 231) (3 downto 2);
                           bin(3 downto 2) <=  TurtokbackString(pixelY - 345, pixelX - 231) (1 downto 0);
              elsif(t1p1(3 downto 0) = "0011") then 
                           rin(3 downto 2) <=  BisaflorbackString(pixelY - 345, pixelX - 231) (5 downto 4);
                           gin(3 downto 2) <=  BisaflorbackString(pixelY - 345, pixelX - 231) (3 downto 2);
                           bin(3 downto 2) <=  BisaflorbackString(pixelY - 345, pixelX - 231) (1 downto 0);
              elsif(t1p1(3 downto 0) = "0100") then
                           rin(3 downto 2) <=  KokoweibackString(pixelY - 345, pixelX - 231) (5 downto 4);
                           gin(3 downto 2) <=  KokoweibackString(pixelY - 345, pixelX - 231) (3 downto 2);
                           bin(3 downto 2) <=  KokoweibackString(pixelY - 345, pixelX - 231) (1 downto 0);
              elsif(t1p1(3 downto 0) = "0101") then 
                           rin(3 downto 2) <=  SarzeniabackString(pixelY - 345, pixelX - 231) (5 downto 4);
                           gin(3 downto 2) <=  SarzeniabackString(pixelY - 345, pixelX - 231) (3 downto 2);
                           bin(3 downto 2) <=  SarzeniabackString(pixelY - 345, pixelX - 231) (1 downto 0);
              elsif(t1p1(3 downto 0) = "0110") then 
                           rin(3 downto 2) <=  GlurakbackString(pixelY - 345, pixelX - 231) (5 downto 4);
                           gin(3 downto 2) <=  GlurakbackString(pixelY - 345, pixelX - 231) (3 downto 2);
                           bin(3 downto 2) <=  GlurakbackString(pixelY - 345, pixelX - 231) (1 downto 0);
              elsif(t1p1(3 downto 0) = "0111") then 
                           rin(3 downto 2) <=  MagmarbackString(pixelY - 345, pixelX - 231) (5 downto 4);
                           gin(3 downto 2) <=  MagmarbackString(pixelY - 345, pixelX - 231) (3 downto 2);
                           bin(3 downto 2) <=  MagmarbackString(pixelY - 345, pixelX - 231) (1 downto 0);
              elsif(t1p1(3 downto 0) = "1000") then 
                           rin(3 downto 2) <=  GallopabackString(pixelY - 345, pixelX - 231) (5 downto 4);
                           gin(3 downto 2) <=  GallopabackString(pixelY - 345, pixelX - 231) (3 downto 2);
                           bin(3 downto 2) <=  GallopabackString(pixelY - 345, pixelX - 231) (1 downto 0);  
              end if;   
             
            
          --T1P2
          elsif(pixelY > 344 and pixelY < 401 and PixelX > 89 and PixelX < 145 and PAliveStatus(1) = '1') then
              if(T1P2(3 downto 0) = "0000") then
                            rin(3 downto 2) <=  AustossFrontString(pixelY - 345, pixelX - 90) (5 downto 4);
                            gin(3 downto 2) <=  AustossFrontString(pixelY - 345, pixelX - 90) (3 downto 2);
                            bin(3 downto 2) <=  AustossFrontString(pixelY - 345, pixelX - 90) (1 downto 0); 
              elsif(T1P2(3 downto 0) = "0001") then
                            rin(3 downto 2) <=  GaradosFrontString(pixelY - 345, pixelX - 90) (5 downto 4);
                            gin(3 downto 2) <=  GaradosFrontString(pixelY - 345, pixelX - 90) (3 downto 2);
                            bin(3 downto 2) <=  GaradosFrontString(pixelY - 345, pixelX - 90) (1 downto 0);
              elsif(T1P2(3 downto 0) = "0010") then 
                            rin(3 downto 2) <=  TurtokFrontString(pixelY - 345, pixelX - 90) (5 downto 4);
                            gin(3 downto 2) <=  TurtokFrontString(pixelY - 345, pixelX - 90) (3 downto 2);
                            bin(3 downto 2) <=  TurtokFrontString(pixelY - 345, pixelX - 90) (1 downto 0);
              elsif(T1P2(3 downto 0) = "0011") then 
                            rin(3 downto 2) <=  BisaflorFrontString(pixelY - 345, pixelX - 90) (5 downto 4);
                            gin(3 downto 2) <=  BisaflorFrontString(pixelY - 345, pixelX - 90) (3 downto 2);
                            bin(3 downto 2) <=  BisaflorFrontString(pixelY - 345, pixelX - 90) (1 downto 0);
              elsif(T1P2(3 downto 0) = "0100") then
                            rin(3 downto 2) <=  KokoweiFrontString(pixelY - 345, pixelX - 90) (5 downto 4);
                            gin(3 downto 2) <=  KokoweiFrontString(pixelY - 345, pixelX - 90) (3 downto 2);
                            bin(3 downto 2) <=  KokoweiFrontString(pixelY - 345, pixelX - 90) (1 downto 0);
              elsif(T1P2(3 downto 0) = "0101") then 
                            rin(3 downto 2) <=  SarzeniaFrontString(pixelY - 345, pixelX - 90) (5 downto 4);
                            gin(3 downto 2) <=  SarzeniaFrontString(pixelY - 345, pixelX - 90) (3 downto 2);
                            bin(3 downto 2) <=  SarzeniaFrontString(pixelY - 345, pixelX - 90) (1 downto 0);
              elsif(T1P2(3 downto 0) = "0110") then 
                            rin(3 downto 2) <=  GlurakFrontString(pixelY - 345, pixelX - 90) (5 downto 4);
                            gin(3 downto 2) <=  GlurakFrontString(pixelY - 345, pixelX - 90) (3 downto 2);
                            bin(3 downto 2) <=  GlurakFrontString(pixelY - 345, pixelX - 90) (1 downto 0);
              elsif(T1P2(3 downto 0) = "0111") then 
                            rin(3 downto 2) <=  MagmarFrontString(pixelY - 345, pixelX - 90) (5 downto 4);
                            gin(3 downto 2) <=  MagmarFrontString(pixelY - 345, pixelX - 90) (3 downto 2);
                            bin(3 downto 2) <=  MagmarFrontString(pixelY - 345, pixelX - 90) (1 downto 0);
              elsif(T1P2(3 downto 0) = "1000") then 
                            rin(3 downto 2) <=  GallopaFrontString(pixelY - 345, pixelX - 90) (5 downto 4);
                            gin(3 downto 2) <=  GallopaFrontString(pixelY - 345, pixelX - 90) (3 downto 2);
                            bin(3 downto 2) <=  GallopaFrontString(pixelY - 345, pixelX - 90) (1 downto 0);          
              end if;
          
              
                      
          --T2P1
          elsif(pixelY > 214 and pixelY < 270 and PixelX > 500 and PixelX < 556 and PAliveStatus(2) = '1') then
              if(T2P1(3 downto 0) = "0000") then 
                            rin(3 downto 2) <=  AustossFrontString(pixelY - 215, pixelX - 501) (5 downto 4);
                            gin(3 downto 2) <=  AustossFrontString(pixelY - 215, pixelX - 501) (3 downto 2);
                            bin(3 downto 2) <=  AustossFrontString(pixelY - 215, pixelX - 501) (1 downto 0);
              elsif(T2P1(3 downto 0) = "0001") then
                            rin(3 downto 2) <=  GaradosFrontString(pixelY - 215, pixelX - 501) (5 downto 4);
                            gin(3 downto 2) <=  GaradosFrontString(pixelY - 215, pixelX - 501) (3 downto 2);
                            bin(3 downto 2) <=  GaradosFrontString(pixelY - 215, pixelX - 501) (1 downto 0);
              elsif(T2P1(3 downto 0) = "0010") then 
                            rin(3 downto 2) <=  TurtokFrontString(pixelY - 215, pixelX - 501) (5 downto 4);
                            gin(3 downto 2) <=  TurtokFrontString(pixelY - 215, pixelX - 501) (3 downto 2);
                            bin(3 downto 2) <=  TurtokFrontString(pixelY - 215, pixelX - 501) (1 downto 0);
              elsif(T2P1(3 downto 0) = "0011") then 
                            rin(3 downto 2) <=  BisaflorFrontString(pixelY - 215, pixelX - 501) (5 downto 4);
                            gin(3 downto 2) <=  BisaflorFrontString(pixelY - 215, pixelX - 501) (3 downto 2);
                            bin(3 downto 2) <=  BisaflorFrontString(pixelY - 215, pixelX - 501) (1 downto 0);
              elsif(T2P1(3 downto 0) = "0100") then
                            rin(3 downto 2) <=  KokoweiFrontString(pixelY - 215, pixelX - 501) (5 downto 4);
                            gin(3 downto 2) <=  KokoweiFrontString(pixelY - 215, pixelX - 501) (3 downto 2);
                            bin(3 downto 2) <=  KokoweiFrontString(pixelY - 215, pixelX - 501) (1 downto 0);
              elsif(T2P1(3 downto 0) = "0101") then 
                            rin(3 downto 2) <=  SarzeniaFrontString(pixelY - 215, pixelX - 501) (5 downto 4);
                            gin(3 downto 2) <=  SarzeniaFrontString(pixelY - 215, pixelX - 501) (3 downto 2);
                            bin(3 downto 2) <=  SarzeniaFrontString(pixelY - 215, pixelX - 501) (1 downto 0);
              elsif(T2P1(3 downto 0) = "0110") then 
                            rin(3 downto 2) <=  GlurakFrontString(pixelY - 215, pixelX - 501) (5 downto 4);
                            gin(3 downto 2) <=  GlurakFrontString(pixelY - 215, pixelX - 501) (3 downto 2);
                            bin(3 downto 2) <=  GlurakFrontString(pixelY - 215, pixelX - 501) (1 downto 0);
              elsif(T2P1(3 downto 0) = "0111") then 
                            rin(3 downto 2) <=  MagmarFrontString(pixelY - 215, pixelX - 501) (5 downto 4);
                            gin(3 downto 2) <=  MagmarFrontString(pixelY - 215, pixelX - 501) (3 downto 2);
                            bin(3 downto 2) <=  MagmarFrontString(pixelY - 215, pixelX - 501) (1 downto 0);
              elsif(T2P1(3 downto 0) = "1000") then 
                            rin(3 downto 2) <=  GallopaFrontString(pixelY - 215, pixelX - 501) (5 downto 4);
                            gin(3 downto 2) <=  GallopaFrontString(pixelY - 215, pixelX - 501) (3 downto 2);
                            bin(3 downto 2) <=  GallopaFrontString(pixelY - 215, pixelX - 501) (1 downto 0);         
              end if;
         
                      
          --T2P2
          elsif(pixelY > 214 and pixelY < 270 and PixelX > 660 and PixelX < 716 and PAliveStatus(3) = '1') then
              if(T2P2(3 downto 0) = "0000") then 
                            rin(3 downto 2) <=  AustossFrontString(pixelY - 215, pixelX - 661) (5 downto 4);
                            gin(3 downto 2) <=  AustossFrontString(pixelY - 215, pixelX - 661) (3 downto 2);
                            bin(3 downto 2) <=  AustossFrontString(pixelY - 215, pixelX - 661) (1 downto 0);
              elsif(T2P2(3 downto 0) = "0001") then
                            rin(3 downto 2) <=  GaradosFrontString(pixelY - 215, pixelX - 661) (5 downto 4);
                            gin(3 downto 2) <=  GaradosFrontString(pixelY - 215, pixelX - 661) (3 downto 2);
                            bin(3 downto 2) <=  GaradosFrontString(pixelY - 215, pixelX - 661) (1 downto 0);
              elsif(T2P2(3 downto 0) = "0010") then 
                            rin(3 downto 2) <=  TurtokFrontString(pixelY - 215, pixelX - 661) (5 downto 4);
                            gin(3 downto 2) <=  TurtokFrontString(pixelY - 215, pixelX - 661) (3 downto 2);
                            bin(3 downto 2) <=  TurtokFrontString(pixelY - 215, pixelX - 661) (1 downto 0);
              elsif(T2P2(3 downto 0) = "0011") then 
                            rin(3 downto 2) <=  BisaflorFrontString(pixelY - 215, pixelX - 661) (5 downto 4);
                            gin(3 downto 2) <=  BisaflorFrontString(pixelY - 215, pixelX - 661) (3 downto 2);
                            bin(3 downto 2) <=  BisaflorFrontString(pixelY - 215, pixelX - 661) (1 downto 0);
              elsif(T2P2(3 downto 0) = "0100") then
                            rin(3 downto 2) <=  KokoweiFrontString(pixelY - 215, pixelX - 661) (5 downto 4);
                            gin(3 downto 2) <=  KokoweiFrontString(pixelY - 215, pixelX - 661) (3 downto 2);
                            bin(3 downto 2) <=  KokoweiFrontString(pixelY - 215, pixelX - 661) (1 downto 0);
              elsif(T2P2(3 downto 0) = "0101") then 
                            rin(3 downto 2) <=  SarzeniaFrontString(pixelY - 215, pixelX - 661) (5 downto 4);
                            gin(3 downto 2) <=  SarzeniaFrontString(pixelY - 215, pixelX - 661) (3 downto 2);
                            bin(3 downto 2) <=  SarzeniaFrontString(pixelY - 215, pixelX - 661) (1 downto 0);
              elsif(T2P2(3 downto 0) = "0110") then 
                            rin(3 downto 2) <=  GlurakFrontString(pixelY - 215, pixelX - 661) (5 downto 4);
                            gin(3 downto 2) <=  GlurakFrontString(pixelY - 215, pixelX - 661) (3 downto 2);
                            bin(3 downto 2) <=  GlurakFrontString(pixelY - 215, pixelX - 661) (1 downto 0);
              elsif(T2P2(3 downto 0) = "0111") then 
                            rin(3 downto 2) <=  MagmarFrontString(pixelY - 215, pixelX - 661) (5 downto 4);
                            gin(3 downto 2) <=  MagmarFrontString(pixelY - 215, pixelX - 661) (3 downto 2);
                            bin(3 downto 2) <=  MagmarFrontString(pixelY - 215, pixelX - 661) (1 downto 0);
              elsif(T2P2(3 downto 0) = "1000") then 
                            rin(3 downto 2) <=  GallopaFrontString(pixelY - 215, pixelX - 661) (5 downto 4);
                            gin(3 downto 2) <=  GallopaFrontString(pixelY - 215, pixelX - 661) (3 downto 2);
                            bin(3 downto 2) <=  GallopaFrontString(pixelY - 215, pixelX - 661) (1 downto 0);   
              end if;            
          end if;
          
          
          
          
          --First Attack Determiner
          if (Bmenu = "000") then
          
          --First Choses
          elsif (Bmenu = "001") then
          
          --Team
            if(pixelX > 298 and pixelX < 386 and pixelY > 100 and pixelY < 134) then
                  if(teamstring(pixely-101, pixelx-299) = '0') then
                  rin <= "0000";
                  gin <= "0000";
                  bin <= "0000";
                  else
                  rin <= "1111";
                  gin <= "1111";
                  bin <= "1111";
                  end if;
              end if;
              
             --1
            if(pixelx > 392 and pixelx < 408 and pixely > 100 and pixely < 134) then
              if(onestring(pixely -101, pixelx-393) = '0') then
                  rin <= "0000";
                  gin <= "0000";
                  bin <= "0000";
              else
                  rin <= "1111";
                  gin <= "1111";
                  bin <= "1111";
              end if;
             end if;
             
             --plays  
            if(pixelx > 415 and pixelx < 504 and pixely > 100 and pixely < 139) then
               if(playsstring(pixely -101, pixelx-416) = '0') then
                   rin <= "0000";
                   gin <= "0000";
                   bin <= "0000";
               else
                   rin <= "1111";
                   gin <= "1111";
                   bin <= "1111";
               end if;
              end if;
            
            --MegaPunch
            if(pixelY > 446 and pixelY < 475 and PixelX > 410 and PixelX < 547) then
                if(MegaPunchString(PixelY - 447, PixelX - 411) = '0') then
                rin <= "0000";
                gin <= "0000";
                bin <= "0000";
                
                else
                rin <= "1111";
                gin <= "1111";
                bin <= "1111";
                end if;
             end if;
             
             --Surf
                   if( (t1p1(3 downto 0) = "0000") or (t1p1(3 downto 0) = "0001") or (t1p1(3 downto 0) = "0010")) then
                    
                    if(pixelY > 448 and pixelY < 471 and PixelX > 342 and PixelX < 390) then
                         if(SurfString(PixelY - 449, PixelX - 343) = '0') then
                         rin <= "0000";
                         gin <= "0000";
                         bin <= "0000";
                         
                         else
                         rin <= "1111";
                         gin <= "1111";
                         bin <= "1111";
                         end if;
                    end if;
                   --LeafBlade
                   elsif( t1p1(3 downto 0) = "0011" or t1p1(3 downto 0) = "0100" or t1p1(3 downto 0) = "0101") then
                   
                     if(pixelY > 448 and pixelY < 473 and PixelX > 274 and PixelX < 390) then
                         if(LeafBladeString(PixelY - 449, PixelX - 275) = '0') then
                         rin <= "0000";
                         gin <= "0000";
                         bin <= "0000";
                         
                         else
                         rin <= "1111";
                         gin <= "1111";
                         bin <= "1111";
                         end if;
                    end if;
                    
                   --FireBlast
                   elsif( t1p1(3 downto 0) = "0110" or t1p1(3 downto 0) = "0111" or t1p1(3 downto 0) = "1000") then
                   
                     if(pixelY > 443 and pixelY < 473 and PixelX > 293 and PixelX < 390) then
                         if(FireBlastString(PixelY - 444, PixelX - 294) = '0') then
                         rin <= "0000";
                         gin <= "0000";
                         bin <= "0000";
                         
                         else
                         rin <= "1111";
                         gin <= "1111";
                         bin <= "1111";
                         end if;
                    end if;           
                   end if;
            
          
          --Second Choses 
          elsif (Bmenu = "011") then
              --team
              if(pixelX > 298 and pixelX < 386 and pixelY > 100 and pixelY < 134) then
                    if(teamstring(pixely-101, pixelx-299) = '0') then
                    rin <= "0000";
                    gin <= "0000";
                    bin <= "0000";
                    else
                    rin <= "1111";
                    gin <= "1111";
                    bin <= "1111";
                    end if;
                end if;
                
               --2
               if(pixelx > 389 and pixelx < 412 and pixely > 100 and pixely < 134) then
                   if(twostring(pixely -101, pixelx-390) = '0') then
                       rin <= "0000";
                       gin <= "0000";
                       bin <= "0000";
                   else
                       rin <= "1111";
                       gin <= "1111";
                       bin <= "1111";
                   end if;
               end if;
               
               --plays  
               if(pixelx > 415 and pixelx < 504 and pixely > 100 and pixely < 139) then
                  if(playsstring(pixely -101, pixelx-416) = '0') then
                      rin <= "0000";
                      gin <= "0000";
                      bin <= "0000";
                  else
                      rin <= "1111";
                      gin <= "1111";
                      bin <= "1111";
                  end if;
                 end if;
                
                        
              --MegaPunch
              if((pixelY > 446 and pixelY < 475 and PixelX > 410 and PixelX < 547)) then
                  if(MegaPunchString(PixelY - 447, PixelX - 411) = '0') then
                  rin <= "0000";
                  gin <= "0000";
                  bin <= "0000";
                  
                  else
                  rin <= "1111";
                  gin <= "1111";
                  bin <= "1111";
                  end if;
               end if;
               
                --Surf
                                 if( (t2p1(3 downto 0) = "0000") or (t2p1(3 downto 0) = "0001") or (t2p1(3 downto 0) = "0010")) then
                                  
                                  if(pixelY > 448 and pixelY < 471 and PixelX > 342 and PixelX < 390) then
                                       if(SurfString(PixelY - 449, PixelX - 343) = '0') then
                                       rin <= "0000";
                                       gin <= "0000";
                                       bin <= "0000";
                                       
                                       else
                                       rin <= "1111";
                                       gin <= "1111";
                                       bin <= "1111";
                                       end if;
                                  end if;
                                 --LeafBlade
                                 elsif( t2p1(3 downto 0) = "0011" or t2p1(3 downto 0) = "0100" or t2p1(3 downto 0) = "0101") then
                                 
                                   if(pixelY > 448 and pixelY < 473 and PixelX > 274 and PixelX < 390) then
                                       if(LeafBladeString(PixelY - 449, PixelX - 275) = '0') then
                                       rin <= "0000";
                                       gin <= "0000";
                                       bin <= "0000";
                                       
                                       else
                                       rin <= "1111";
                                       gin <= "1111";
                                       bin <= "1111";
                                       end if;
                                  end if;
                                  
                                 --FireBlast
                                 elsif( t2p1(3 downto 0) = "0110" or t2p1(3 downto 0) = "0111" or t2p1(3 downto 0) = "1000") then
                                 
                                   if(pixelY > 443 and pixelY < 473 and PixelX > 293 and PixelX < 390) then
                                       if(FireBlastString(PixelY - 444, PixelX - 294) = '0') then
                                       rin <= "0000";
                                       gin <= "0000";
                                       bin <= "0000";
                                       
                                       else
                                       rin <= "1111";
                                       gin <= "1111";
                                       bin <= "1111";
                                       end if;
                                  end if;           
                                 end if;
               
          --Damage Screen
          elsif (Bmenu = "100" or Bmenu = "010") then
                
                if(Bmenu= "100" and angriff /= "111") then
                    if (pixelY > 309 and pixelY < 313 and pixelX > 270 +hp1 and pixelX < 270 + hp1 + rot) then
                          rin <= "1111";
                          gin <= "0000";
                          bin <= "0000";
                    end if;
                    
                    --Normale
                    if (pixelY > 363 and pixelY < 380 and pixelX > 248 and pixelX < 268 and  angriff = "000") then
                        if(normaleString(pixely - 364, pixelX - 249) /= "000000") then
                          rin(3 downto 2) <= normaleString(pixely - 364, pixelX - 249)(5 downto 4);
                          gin(3 downto 2) <= normaleString(pixely - 364, pixelX - 249)(3 downto 2);
                          bin(3 downto 2) <= normaleString(pixely - 364, pixelX - 249)(1 downto 0);
                        end if;
                    --Wasser
                    elsif (pixelY > 356 and pixelY < 401 and pixelX > 248 and pixelX < 268 and  angriff = "001") then
                    if(wasserString(pixely - 357, pixelX - 249) /= "000000") then
                          rin(3 downto 2) <= wasserString(pixely - 357, pixelX - 249)(5 downto 4);
                          gin(3 downto 2) <= wasserString(pixely - 357, pixelX - 249)(3 downto 2);
                          bin(3 downto 2) <= wasserString(pixely - 357, pixelX - 249)(1 downto 0);
                          end if;
                    --Feuer
                    elsif (pixelY > 389 and pixelY < 401 and pixelX > 245 and pixelX < 279 and  angriff = "011") then
                          if(feuerString(pixely - 390, pixelX - 246) /= "000000") then
                          rin(3 downto 2) <= feuerString(pixely - 414, pixelX - 246)(5 downto 4);
                          gin(3 downto 2) <= feuerString(pixely - 414, pixelX - 246)(3 downto 2);
                          bin(3 downto 2) <= feuerString(pixely - 414, pixelX - 246)(1 downto 0);
                          end if;
                    --Pflanze
                    elsif (pixelY > 361 and pixelY < 384 and pixelX > 245 and pixelX < 272 and  angriff = "010") then
                          if(pflanzeString(pixely - 362, pixelX - 246) /= "000000") then
                          rin(3 downto 2) <= pflanzeString(pixely - 362, pixelX - 246)(5 downto 4);
                          gin(3 downto 2) <= pflanzeString(pixely - 362, pixelX - 246)(3 downto 2);
                          bin(3 downto 2) <= pflanzeString(pixely - 362, pixelX - 246)(1 downto 0);
                          end if;
                    end if;
                else
                    if (pixelY > 179 and pixelY < 183 and pixelX > 540 +hp2 and pixelX < 540 +hp2 + rot and angriff /= "111") then
                        rin <= "1111";
                        gin <= "0000";
                        bin <= "0000";
                    end if;   
                    
                    --Normale
                    if (pixelY > 233 and pixelY < 250 and pixelX > 518 and pixelX < 538 and  angriff = "000") then
                        if(normaleString(pixely - 234, pixelX - 519) /= "000000") then
                          rin(3 downto 2) <= normaleString(pixely - 234, pixelX - 519)(5 downto 4);
                          gin(3 downto 2) <= normaleString(pixely - 234, pixelX - 519)(3 downto 2);
                          bin(3 downto 2) <= normaleString(pixely - 234, pixelX - 519)(1 downto 0);
                        end if;
                    --Wasser
                    elsif (pixelY > 225 and pixelY < 270 and pixelX > 518 and pixelX < 538 and  angriff = "001") then
                    if(wasserString(pixely - 226, pixelX - 519) /= "000000") then
                          rin(3 downto 2) <= wasserString(pixely - 226, pixelX - 519)(5 downto 4);
                          gin(3 downto 2) <= wasserString(pixely - 226, pixelX - 519)(3 downto 2);
                          bin(3 downto 2) <= wasserString(pixely - 226, pixelX - 519)(1 downto 0);
                          end if;
                    --Feuer
                    elsif (pixelY > 258 and pixelY < 270 and pixelX > 515 and pixelX < 549 and  angriff = "011") then
                          if(feuerString(pixely - 259, pixelX - 516) /= "000000") then
                          rin(3 downto 2) <= feuerString(pixely - 284, pixelX - 516)(5 downto 4);
                          gin(3 downto 2) <= feuerString(pixely - 284, pixelX - 516)(3 downto 2);
                          bin(3 downto 2) <= feuerString(pixely - 284, pixelX - 516)(1 downto 0);
                          end if;
                    --Pflanze
                    elsif (pixelY > 231 and pixelY < 254 and pixelX > 515 and pixelX < 542 and  angriff = "010") then
                          if(pflanzeString(pixely - 232, pixelX - 519) /= "000000") then
                          rin(3 downto 2) <= pflanzeString(pixely - 232, pixelX - 516)(5 downto 4);
                          gin(3 downto 2) <= pflanzeString(pixely - 232, pixelX - 516)(3 downto 2);
                          bin(3 downto 2) <= pflanzeString(pixely - 232, pixelX - 516)(1 downto 0);
                          end if;
                    end if;
                end if; 
                  
                --Surf
                if(angriff = "001") then
                  if (PixelY > 420 and PixelY < 443 and PixelX > 170 and PixelX < 218 ) then
                       if(SurfString(PixelY - 421, PixelX - 171) = '0') then
                       rin <= "0000";
                       gin <= "0000";
                       bin <= "0000";
                       
                       else
                       rin <= "1111";
                       gin <= "1111";
                       bin <= "1111";
                       end if;
                  end if;
                
                --Leaf Blade
                elsif(angriff = "010") then
                  if (PixelY > 420 and PixelY < 445 and PixelX > 170 and PixelX < 286 ) then
                       if(LeafBladeString(PixelY - 421, PixelX - 171) = '0') then
                       rin <= "0000";
                       gin <= "0000";
                       bin <= "0000";
                       
                       else
                       rin <= "1111";
                       gin <= "1111";
                       bin <= "1111";
                       end if;
                  end if;
                --Fire Blast
                elsif(angriff = "011") then
                  if (PixelY > 420 and PixelY < 445 and PixelX > 170 and PixelX < 267 ) then
                       if(FireBlastString(PixelY - 421, PixelX - 171) = '0') then
                       rin <= "0000";
                       gin <= "0000";
                       bin <= "0000";
                       
                       else
                       rin <= "1111";
                       gin <= "1111";
                       bin <= "1111";
                       end if;
                  end if;
                end if;  
                  
                  --MegaPunch
                if (angriff = "000") then
                  if (PixelY > 420 and PixelY < 449 and PixelX > 170 and PixelX < 307 ) then
                       if(MegaPunchString(PixelY - 421, PixelX - 171) = '0') then
                       rin <= "0000";
                       gin <= "0000";
                       bin <= "0000";
                       
                       else
                       rin <= "1111";
                       gin <= "1111";
                       bin <= "1111";
                       end if;
                    end if;  
                  
                 elsif(ddamage = '0' and angriff /= "111") then
                    --not
                    if(PixelY > 455 and PixelY < 472 and PixelX > 170 and PixelX < 207) then
                        if(NotString(PixelY - 456, PixelX - 171) = '0') then
                        rin <= "0000";
                        gin <= "0000";
                        bin <= "0000";
                        
                        else
                        rin <= "1111";
                        gin <= "1111";
                        bin <= "1111";
                        end if;
                      end if;
                      
                      --very effective
                      if(PixelY > 455 and PixelY < 477 and PixelX > 210 and PixelX < 366) then
                        if(VeryEffectiveString(PixelY - 456, PixelX - 211) = '0') then
                        rin <= "0000";
                        gin <= "0000";
                        bin <= "0000";
                        
                        else
                        rin <= "1111";
                        gin <= "1111";
                        bin <= "1111";
                        end if; 
                      end if;  
                 
                  
                  
                elsif(ddamage = '1' and angriff /= "111") then
                --very effective
                  if(PixelY > 455 and PixelY < 477 and PixelX > 170 and PixelX < 326) then
                    if(VeryEffectiveString(PixelY - 456, PixelX - 171) = '0') then
                    rin <= "0000";
                    gin <= "0000";
                    bin <= "0000";
                    
                    else
                    rin <= "1111";
                    gin <= "1111";
                    bin <= "1111";
                    end if; 
                  end if; 
                  
               end if;
          end if;
     
     --Winner
     elsif (menu = "101") then
     --Team
        if(pixelX > 298 and pixelX < 386 and pixelY > 200 and pixelY < 234) then
            if(teamstring(pixely-201, pixelx-299) = '0') then
            rin <= "0000";
            gin <= "0000";
            bin <= "0000";
            else
            rin <= "1111";
            gin <= "1111";
            bin <= "1111";
            end if;
        end if;
        
        --Wins
        if(pixelX > 415 and pixelX < 516 and pixelY > 200 and pixelY < 234) then
            if(winsstring(pixely-201, pixelx-299) = '0') then
            rin <= "0000";
            gin <= "0000";
            bin <= "0000";
            else
            rin <= "1111";
            gin <= "1111";
            bin <= "1111";
            end if;
        end if;
        
        --1 or 2
        if(winner = '0') then
           if(pixelx > 392 and pixelx < 408 and pixely > 200 and pixely < 234) then
            if(onestring(pixely -201, pixelx-393) = '0') then
                rin <= "0000";
                gin <= "0000";
                bin <= "0000";
            else
                rin <= "1111";
                gin <= "1111";
                bin <= "1111";
            end if;
           end if;
         else
            if(pixelx > 389 and pixelx < 412 and pixely > 200 and pixely < 234) then
                if(twostring(pixely -201, pixelx-390) = '0') then
                    rin <= "0000";
                    gin <= "0000";
                    bin <= "0000";
                else
                    rin <= "1111";
                    gin <= "1111";
                    bin <= "1111";
                end if;
            end if;            
         end if;
     end if;
end if;         
end process;



end Behavioral;
